* NGSPICE file created from FC_top.ext - technology: gf180mcuD

.subckt FC_top VP VN VOUT IREF AVSS AVDD
X0 AVDD.t1280 AVDD.t1279 AVDD.t1280 AVDD.t178 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1 AVSS.t282 AVSS.t281 AVSS.t282 AVSS.t43 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2 AVDD.t1376 a_5396_n6451.t67 a_5396_8177.t87 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3 a_n11737_n15980.t23 IREF.t44 AVDD.t1640 AVDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4 AVDD.t1641 IREF.t45 a_n13990_8177.t273 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5 a_5396_8177.t174 a_n11317_n20927.t1 a_5396_n6451.t16 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6 AVDD.t1278 AVDD.t1277 AVDD.t1278 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X7 a_5396_8177.t86 a_5396_n6451.t68 AVDD.t1377 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X8 AVDD.t1276 AVDD.t1275 AVDD.t1276 AVDD.t373 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X9 AVDD.t1642 IREF.t46 a_n13990_8177.t272 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X10 AVDD.t1643 IREF.t47 a_n13990_8177.t271 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X11 a_n13990_8177.t1 VP.t0 a_n13990_n6451.t141 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X12 a_n13990_n5465.t112 VN.t0 a_n13990_8177.t303 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X13 VOUT.t87 a_n11317_n20927.t1 a_5396_9163.t137 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X14 a_n13990_n5465.t111 VN.t1 a_n13990_8177.t304 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X15 AVDD.t1644 IREF.t48 a_n13990_8177.t270 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X16 a_n13990_n6451.t140 VP.t1 a_n13990_8177.t0 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X17 a_5396_8177.t173 a_n11317_n20927.t1 a_5396_n6451.t16 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X18 AVDD.t1274 AVDD.t1273 AVDD.t1274 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X19 a_n13990_8177.t92 VP.t2 a_n13990_n6451.t139 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X20 a_n13990_n5465.t110 VN.t2 a_n13990_8177.t305 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X21 AVDD.t1645 IREF.t49 a_n13990_8177.t269 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X22 AVDD.t1272 AVDD.t1271 AVDD.t1272 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X23 AVDD.t1270 AVDD.t1269 AVDD.t1270 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X24 a_n11737_n15980.t22 IREF.t50 AVDD.t1646 AVDD.t39 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X25 a_n13990_8177.t268 IREF.t51 AVDD.t1647 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X26 a_n13990_8177.t267 IREF.t52 AVDD.t1648 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X27 AVDD.t1268 AVDD.t1267 AVDD.t1268 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X28 AVDD.t1266 AVDD.t1265 AVDD.t1266 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X29 AVSS.t280 AVSS.t279 AVSS.t280 AVSS.t74 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X30 AVDD.t1378 a_5396_n6451.t69 a_5396_9163.t87 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X31 AVDD.t1264 AVDD.t1263 AVDD.t1264 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X32 a_5396_9163.t86 a_5396_n6451.t70 AVDD.t1528 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X33 a_5396_9163.t85 a_5396_n6451.t71 AVDD.t1529 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X34 AVDD.t1262 AVDD.t1261 AVDD.t1262 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X35 AVDD.t1604 IREF.t42 IREF.t43 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X36 AVDD.t1260 AVDD.t1259 AVDD.t1260 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X37 AVDD.t1530 a_5396_n6451.t72 a_5396_9163.t84 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X38 AVDD.t1649 IREF.t53 a_n13990_8177.t266 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X39 VOUT.t86 a_n11317_n20927.t1 a_5396_9163.t136 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X40 AVDD.t1258 AVDD.t1257 AVDD.t1258 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X41 a_n13990_n6451.t138 VP.t3 a_n13990_8177.t47 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X42 a_5396_n6451.t20 a_n11317_n20927.t1 a_5396_8177.t172 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X43 a_n11737_n15980.t21 IREF.t54 AVDD.t1650 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X44 AVSS.t278 AVSS.t277 AVSS.t278 AVSS.t1 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X45 AVSS.t276 AVSS.t275 AVSS.t276 AVSS.t49 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X46 AVDD.t1651 IREF.t55 a_n11737_n14973.t29 AVDD.t810 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X47 AVDD.t1256 AVDD.t1255 AVDD.t1256 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X48 a_n13990_n5465.t109 VN.t3 a_n13990_8177.t306 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X49 AVDD.t1254 AVDD.t1253 AVDD.t1254 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X50 AVDD.t1252 AVDD.t1251 AVDD.t1252 AVDD.t875 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X51 AVSS.t338 a_n11737_n14973.t30 a_n13990_n5465.t23 AVSS.t82 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X52 AVDD.t1250 AVDD.t1249 AVDD.t1250 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X53 AVDD.t1248 AVDD.t1247 AVDD.t1248 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X54 a_n13990_n5465.t24 a_n11737_n14973.t31 AVSS.t339 AVSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X55 a_5396_8177.t171 a_n11317_n20927.t1 a_5396_n6451.t19 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X56 AVSS.t274 AVSS.t273 AVSS.t274 AVSS.t55 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X57 a_5396_8177.t85 a_5396_n6451.t73 AVDD.t1531 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X58 a_n1533_n15598# a_n11317_n20927.t3 a_n2101_n15598# AVDD.t394 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X59 a_5396_8177.t84 a_5396_n6451.t74 AVDD.t1532 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X60 AVDD.t1533 a_5396_n6451.t75 a_5396_9163.t83 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X61 a_n13990_8177.t265 IREF.t56 AVDD.t1652 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X62 AVDD.t1246 AVDD.t1245 AVDD.t1246 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X63 VOUT.t85 a_n11317_n20927.t1 a_5396_9163.t143 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X64 a_5396_8177.t170 a_n11317_n20927.t1 a_5396_n6451.t18 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X65 AVDD.t1244 AVDD.t1243 AVDD.t1244 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X66 a_n13990_n5465.t15 a_n11737_n14973.t32 AVSS.t321 AVSS.t158 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X67 AVDD.t1653 IREF.t57 a_n11737_n15980.t20 AVDD.t810 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X68 a_n13990_n5465.t16 a_n11737_n14973.t33 AVSS.t322 AVSS.t155 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X69 a_n13990_n5465.t108 VN.t4 a_n13990_8177.t317 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X70 AVDD.t1242 AVDD.t1241 AVDD.t1242 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X71 a_n13990_8177.t264 IREF.t58 AVDD.t1654 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X72 AVDD.t1655 IREF.t59 a_n13990_8177.t263 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X73 a_5396_n6451.t17 a_n11317_n20927.t1 a_5396_8177.t169 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X74 a_5396_n6451.t16 a_n11317_n20927.t1 a_5396_8177.t168 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X75 a_5396_9163.t142 a_n11317_n20927.t1 VOUT.t84 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X76 AVSS.t272 AVSS.t271 AVSS.t272 AVSS.t25 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X77 a_n13990_n5465.t17 a_n11737_n14973.t34 AVSS.t323 AVSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X78 a_n13990_n6451.t48 a_n11737_n15980.t24 a_5396_n6451.t65 AVSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X79 a_n11317_n20927.t1 a_n11737_n14973.t35 AVSS.t324 AVSS.t31 nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X80 AVDD.t1240 AVDD.t1239 AVDD.t1240 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X81 VOUT.t83 a_n11317_n20927.t1 a_5396_9163.t157 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X82 a_n13990_8177.t279 VP.t4 a_n13990_n6451.t137 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X83 AVDD.t1238 AVDD.t1237 AVDD.t1238 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X84 AVDD.t1236 AVDD.t1235 AVDD.t1236 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X85 a_5396_n6451.t15 a_n11317_n20927.t1 a_5396_8177.t167 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X86 AVDD.t1534 a_5396_n6451.t76 a_5396_8177.t83 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X87 a_n13990_8177.t262 IREF.t60 AVDD.t1656 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X88 a_5396_9163.t156 a_n11317_n20927.t1 VOUT.t82 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X89 AVDD.t1234 AVDD.t1233 AVDD.t1234 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X90 a_5396_n6451.t16 a_n11317_n20927.t1 a_5396_8177.t166 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X91 AVDD.t1232 AVDD.t1231 AVDD.t1232 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X92 a_5396_8177.t82 a_5396_n6451.t77 AVDD.t1535 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X93 AVDD.t1536 a_5396_n6451.t78 a_5396_9163.t82 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X94 AVDD.t1230 AVDD.t1229 AVDD.t1230 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X95 AVDD.t1537 a_5396_n6451.t79 a_5396_9163.t81 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X96 a_n13990_8177.t280 VP.t5 a_n13990_n6451.t136 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X97 AVDD.t1228 AVDD.t1227 AVDD.t1228 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X98 AVDD.t1226 AVDD.t1225 AVDD.t1226 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X99 AVDD.t1580 IREF.t61 a_n13990_8177.t261 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X100 AVDD.t1581 IREF.t62 a_n13990_8177.t260 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X101 AVDD.t1224 AVDD.t1223 AVDD.t1224 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X102 a_n13990_8177.t259 IREF.t63 AVDD.t1582 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X103 a_5396_9163.t80 a_5396_n6451.t80 AVDD.t1538 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X104 a_5396_n6451.t24 a_n11317_n20927.t1 a_5396_8177.t165 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X105 a_5396_8177.t164 a_n11317_n20927.t1 a_5396_n6451.t49 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X106 AVDD.t1222 AVDD.t1221 AVDD.t1222 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X107 AVSS.t270 AVSS.t269 AVSS.t270 AVSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X108 AVDD.t1220 AVDD.t1219 AVDD.t1220 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X109 AVDD.t1218 AVDD.t1217 AVDD.t1218 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X110 a_n1533_n16323# a_n11317_n20927.t1 a_n2101_n16323# AVDD.t394 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X111 a_n13990_8177.t258 IREF.t64 AVDD.t1583 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X112 AVSS.t268 AVSS.t267 AVSS.t268 AVSS.t235 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X113 VOUT.t81 a_n11317_n20927.t1 a_5396_9163.t147 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X114 AVDD.t1216 AVDD.t1215 AVDD.t1216 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X115 a_5396_9163.t79 a_5396_n6451.t81 AVDD.t1539 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X116 AVDD.t1214 AVDD.t1213 AVDD.t1214 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X117 AVDD.t1584 IREF.t65 a_n13990_8177.t257 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X118 AVDD.t1212 AVDD.t1211 AVDD.t1212 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X119 AVDD.t1210 AVDD.t1209 AVDD.t1210 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X120 AVDD.t1208 AVDD.t1207 AVDD.t1208 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X121 IREF.t41 IREF.t40 AVDD.t1603 AVDD.t480 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X122 a_n11737_n14973.t28 IREF.t66 AVDD.t1585 AVDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X123 AVDD.t1206 AVDD.t1205 AVDD.t1206 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X124 a_n13990_n6451.t135 VP.t6 a_n13990_8177.t281 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X125 AVDD.t1204 AVDD.t1203 AVDD.t1204 AVDD.t810 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X126 AVDD.t1202 AVDD.t1201 AVDD.t1202 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X127 AVDD.t1586 IREF.t67 a_n13990_8177.t256 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X128 AVDD.t1587 IREF.t68 a_n11737_n15980.t19 AVDD.t638 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X129 AVDD.t1588 IREF.t69 a_n13990_8177.t255 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X130 VOUT.t80 a_n11317_n20927.t1 a_5396_9163.t146 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X131 a_5396_9163.t78 a_5396_n6451.t82 AVDD.t1540 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X132 AVDD.t1200 AVDD.t1199 AVDD.t1200 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X133 AVDD.t1589 IREF.t70 a_n13990_8177.t254 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X134 AVDD.t1541 a_5396_n6451.t83 a_5396_8177.t81 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X135 AVDD.t1590 IREF.t71 a_n13990_8177.t253 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X136 a_n13990_8177.t252 IREF.t72 AVDD.t1591 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X137 AVDD.t1592 IREF.t73 a_n13990_8177.t251 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X138 a_n13990_n6451.t11 a_n11737_n14973.t36 AVSS.t299 AVSS.t144 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X139 a_n2101_n15598# a_n11317_n20927.t3 a_n2631_n16323# AVDD.t328 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X140 a_n13990_n6451.t12 a_n11737_n14973.t37 AVSS.t300 AVSS.t141 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X141 AVDD.t1198 AVDD.t1197 AVDD.t1198 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X142 AVDD.t1196 AVDD.t1195 AVDD.t1196 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X143 AVDD.t1194 AVDD.t1193 AVDD.t1194 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X144 AVDD.t1192 AVDD.t1191 AVDD.t1192 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X145 AVDD.t1593 IREF.t74 a_n13990_8177.t250 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X146 AVDD.t1190 AVDD.t1189 AVDD.t1190 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X147 AVDD.t1188 AVDD.t1187 AVDD.t1188 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X148 AVDD.t1186 AVDD.t1185 AVDD.t1186 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X149 AVDD.t1542 a_5396_n6451.t84 a_5396_8177.t80 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X150 a_n13990_8177.t249 IREF.t75 AVDD.t1594 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X151 a_5396_n6451.t48 a_n11317_n20927.t1 a_5396_8177.t163 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X152 AVDD.t1184 AVDD.t1183 AVDD.t1184 AVDD.t264 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X153 AVDD.t1182 AVDD.t1181 AVDD.t1182 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X154 a_n13990_n5465.t126 a_n11737_n15980.t25 VOUT.t105 AVSS.t88 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X155 a_n13990_n5465.t125 a_n11737_n15980.t26 VOUT.t104 AVSS.t85 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X156 AVDD.t1595 IREF.t76 a_n11737_n15980.t18 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X157 a_n13990_8177.t248 IREF.t77 AVDD.t1596 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X158 a_5396_8177.t162 a_n11317_n20927.t1 a_5396_n6451.t47 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X159 VOUT.t79 a_n11317_n20927.t1 a_5396_9163.t101 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X160 a_n13990_n5465.t107 VN.t5 a_n13990_8177.t318 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X161 AVDD.t1180 AVDD.t1179 AVDD.t1180 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X162 IREF.t39 IREF.t38 AVDD.t1602 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X163 AVDD.t1178 AVDD.t1177 AVDD.t1178 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X164 a_n13990_8177.t247 IREF.t78 AVDD.t1674 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X165 AVDD.t1176 AVDD.t1175 AVDD.t1176 AVDD.t156 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X166 AVSS.t266 AVSS.t265 AVSS.t266 AVSS.t28 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X167 AVDD.t1675 IREF.t79 a_n13990_8177.t246 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X168 AVDD.t1543 a_5396_n6451.t85 a_5396_8177.t79 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X169 a_5396_8177.t78 a_5396_n6451.t86 AVDD.t1544 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X170 AVDD.t1174 AVDD.t1173 AVDD.t1174 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X171 a_n13990_8177.t282 VP.t7 a_n13990_n6451.t134 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X172 AVDD.t1545 a_5396_n6451.t87 a_5396_9163.t77 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X173 AVDD.t1546 a_5396_n6451.t88 a_5396_8177.t77 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X174 AVDD.t1172 AVDD.t1171 AVDD.t1172 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X175 AVDD.t1170 AVDD.t1169 AVDD.t1170 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X176 a_5396_8177.t161 a_n11317_n20927.t1 a_5396_n6451.t47 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X177 a_n13990_n5465.t106 VN.t6 a_n13990_8177.t319 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X178 VOUT.t78 a_n11317_n20927.t1 a_5396_9163.t100 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X179 AVDD.t1676 IREF.t80 a_n11737_n14973.t27 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X180 AVSS.t264 AVSS.t263 AVSS.t264 AVSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X181 AVSS.t262 AVSS.t261 AVSS.t262 AVSS.t16 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X182 AVSS.t260 AVSS.t259 AVSS.t260 AVSS.t19 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X183 AVDD.t1168 AVDD.t1167 AVDD.t1168 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X184 a_5396_9163.t173 a_n11317_n20927.t1 VOUT.t77 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X185 AVDD.t1677 IREF.t81 a_n11737_n14973.t26 AVDD.t282 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X186 a_5396_9163.t172 a_n11317_n20927.t1 VOUT.t76 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X187 a_n13990_n6451.t133 VP.t8 a_n13990_8177.t327 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X188 a_n13990_8177.t328 VP.t9 a_n13990_n6451.t132 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X189 a_n2101_n16323# a_n11317_n20927.t1 a_n2631_n16323# AVDD.t328 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X190 a_5396_n6451.t46 a_n11317_n20927.t1 a_5396_8177.t160 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X191 VOUT.t75 a_n11317_n20927.t1 a_5396_9163.t127 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X192 AVDD.t1547 a_5396_n6451.t89 a_5396_8177.t76 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X193 a_5396_9163.t76 a_5396_n6451.t90 AVDD.t1548 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X194 AVSS.t301 a_n11737_n14973.t38 a_n13990_n6451.t13 AVSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X195 a_n6139_n21443# a_n11737_n15980.t27 a_n6661_n21443# AVSS.t178 nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X196 a_5396_9163.t75 a_5396_n6451.t91 AVDD.t1549 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X197 a_n13990_n5465.t130 a_n11737_n15980.t28 VOUT.t103 AVSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X198 AVDD.t1166 AVDD.t1165 AVDD.t1166 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X199 a_5396_8177.t75 a_5396_n6451.t92 AVDD.t1550 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X200 AVDD.t1164 AVDD.t1163 AVDD.t1164 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X201 a_5396_n6451.t45 a_n11317_n20927.t1 a_5396_8177.t159 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X202 AVDD.t1162 AVDD.t1161 AVDD.t1162 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X203 AVDD.t1678 IREF.t82 a_n13990_8177.t245 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X204 AVSS.t302 a_n11737_n14973.t39 a_n13990_n6451.t14 AVSS.t114 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X205 a_5396_9163.t126 a_n11317_n20927.t1 VOUT.t74 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X206 a_n13990_8177.t320 VN.t7 a_n13990_n5465.t105 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X207 AVDD.t1160 AVDD.t1159 AVDD.t1160 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X208 VOUT.t73 a_n11317_n20927.t1 a_5396_9163.t91 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X209 a_n13990_8177.t321 VN.t8 a_n13990_n5465.t104 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X210 AVDD.t1158 AVDD.t1157 AVDD.t1158 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X211 a_n13990_8177.t244 IREF.t83 AVDD.t1679 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X212 AVSS.t258 AVSS.t257 AVSS.t258 AVSS.t222 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X213 VOUT.t72 a_n11317_n20927.t1 a_5396_9163.t90 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X214 AVDD.t1156 AVDD.t1155 AVDD.t1156 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X215 AVDD.t1154 AVDD.t1153 AVDD.t1154 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X216 AVDD.t1152 AVDD.t1151 AVDD.t1152 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X217 AVDD.t1150 AVDD.t1149 AVDD.t1150 AVDD.t13 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X218 a_n13990_8177.t347 VN.t9 a_n13990_n5465.t103 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X219 AVDD.t1551 a_5396_n6451.t93 a_5396_8177.t74 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X220 a_5396_9163.t167 a_n11317_n20927.t1 VOUT.t71 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X221 AVDD.t1148 AVDD.t1147 AVDD.t1148 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X222 AVDD.t1146 AVDD.t1145 AVDD.t1146 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X223 a_n13990_n5465.t102 VN.t10 a_n13990_8177.t348 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X224 a_n13990_8177.t349 VN.t11 a_n13990_n5465.t101 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X225 AVDD.t1144 AVDD.t1143 AVDD.t1144 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X226 VOUT.t70 a_n11317_n20927.t1 a_5396_9163.t166 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X227 a_n1533_n17634# a_n11317_n20927.t1 a_n2101_n17634# AVDD.t394 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X228 a_5396_n6451.t14 a_n11317_n20927.t1 a_5396_8177.t158 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X229 AVDD.t1142 AVDD.t1141 AVDD.t1142 AVDD.t181 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X230 AVSS.t256 AVSS.t255 AVSS.t256 AVSS.t28 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X231 AVDD.t1140 AVDD.t1139 AVDD.t1140 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X232 AVDD.t1138 AVDD.t1137 AVDD.t1138 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X233 AVDD.t1136 AVDD.t1135 AVDD.t1136 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X234 AVSS.t254 AVSS.t253 AVSS.t254 AVSS.t1 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X235 AVSS.t334 a_n11737_n14973.t40 a_n13990_n6451.t25 AVSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X236 AVDD.t1134 AVDD.t1133 AVDD.t1134 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X237 AVDD.t1132 AVDD.t1131 AVDD.t1132 AVDD.t373 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X238 a_5396_n6451.t66 a_n11737_n15980.t29 a_n13990_n6451.t47 AVSS.t67 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X239 a_n13990_8177.t350 VN.t12 a_n13990_n5465.t100 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X240 a_5396_n6451.t0 a_n11737_n15980.t30 a_n13990_n6451.t46 AVSS.t64 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X241 AVDD.t1130 AVDD.t1129 AVDD.t1130 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X242 AVDD.t1680 IREF.t84 a_n13990_8177.t243 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X243 AVDD.t1128 AVDD.t1127 AVDD.t1128 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X244 AVDD.t1126 AVDD.t1125 AVDD.t1126 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X245 AVDD.t1552 a_5396_n6451.t94 a_5396_9163.t74 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X246 AVDD.t1681 IREF.t85 a_n13990_8177.t242 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X247 AVDD.t1124 AVDD.t1123 AVDD.t1124 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X248 AVDD.t1122 AVDD.t1121 AVDD.t1122 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X249 AVDD.t1120 AVDD.t1119 AVDD.t1120 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X250 AVDD.t1118 AVDD.t1117 AVDD.t1118 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X251 AVSS.t252 AVSS.t251 AVSS.t252 AVSS.t55 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X252 AVDD.t1116 AVDD.t1115 AVDD.t1116 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X253 AVDD.t1114 AVDD.t1113 AVDD.t1114 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X254 AVDD.t1682 IREF.t86 a_n13990_8177.t241 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X255 AVDD.t1112 AVDD.t1111 AVDD.t1112 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X256 AVDD.t1601 IREF.t36 IREF.t37 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X257 AVDD.t1600 IREF.t34 IREF.t35 AVDD.t638 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X258 AVSS.t250 AVSS.t249 AVSS.t250 AVSS.t74 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X259 AVDD.t1110 AVDD.t1109 AVDD.t1110 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X260 a_n13990_8177.t240 IREF.t87 AVDD.t1683 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X261 a_n13990_n6451.t131 VP.t10 a_n13990_8177.t329 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X262 AVDD.t1108 AVDD.t1107 AVDD.t1108 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X263 AVDD.t1106 AVDD.t1105 AVDD.t1106 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X264 AVDD.t1104 AVDD.t1103 AVDD.t1104 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X265 AVDD.t1102 AVDD.t1101 AVDD.t1102 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X266 AVDD.t1100 AVDD.t1099 AVDD.t1100 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X267 AVDD.t1098 AVDD.t1097 AVDD.t1098 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X268 AVDD.t1096 AVDD.t1095 AVDD.t1096 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X269 a_n13990_8177.t330 VP.t11 a_n13990_n6451.t130 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X270 a_5396_8177.t73 a_5396_n6451.t95 AVDD.t1553 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X271 AVDD.t1094 AVDD.t1093 AVDD.t1094 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X272 a_n13990_8177.t331 VP.t12 a_n13990_n6451.t129 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X273 AVDD.t1092 AVDD.t1091 AVDD.t1092 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X274 AVDD.t1684 IREF.t88 a_n13990_8177.t239 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X275 a_n11737_n14973.t25 IREF.t89 AVDD.t1685 AVDD.t638 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X276 AVDD.t1090 AVDD.t1089 AVDD.t1090 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X277 AVDD.t1088 AVDD.t1087 AVDD.t1088 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X278 AVDD.t1086 AVDD.t1085 AVDD.t1086 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X279 VOUT.t69 a_n11317_n20927.t1 a_5396_9163.t115 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X280 AVDD.t1686 IREF.t90 a_n13990_8177.t238 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X281 AVSS.t248 AVSS.t247 AVSS.t248 AVSS.t138 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X282 AVDD.t1084 AVDD.t1083 AVDD.t1084 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X283 AVSS.t246 AVSS.t245 AVSS.t246 AVSS.t46 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X284 AVDD.t1687 IREF.t91 a_n13990_8177.t237 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X285 VOUT.t68 a_n11317_n20927.t1 a_5396_9163.t114 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X286 AVDD.t1082 AVDD.t1081 AVDD.t1082 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X287 a_n13990_8177.t236 IREF.t92 AVDD.t1688 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X288 AVDD.t1080 AVDD.t1079 AVDD.t1080 AVDD.t131 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X289 AVDD.t1078 AVDD.t1077 AVDD.t1078 AVDD.t193 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X290 a_5396_n6451.t4 a_n11737_n15980.t31 a_n13990_n6451.t45 AVSS.t88 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X291 AVDD.t1076 AVDD.t1075 AVDD.t1076 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X292 a_5396_n6451.t1 a_n11737_n15980.t32 a_n13990_n6451.t44 AVSS.t85 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X293 AVDD.t1074 AVDD.t1073 AVDD.t1074 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X294 AVDD.t1072 AVDD.t1071 AVDD.t1072 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X295 AVDD.t1070 AVDD.t1069 AVDD.t1070 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X296 AVDD.t1068 AVDD.t1067 AVDD.t1068 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X297 a_n13990_8177.t235 IREF.t93 AVDD.t1689 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X298 a_n13990_n6451.t43 a_n11737_n15980.t33 a_5396_n6451.t1 AVSS.t37 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X299 AVDD.t1066 AVDD.t1065 AVDD.t1066 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X300 AVDD.t1554 a_5396_n6451.t96 a_5396_9163.t73 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X301 AVDD.t1064 AVDD.t1063 AVDD.t1064 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X302 a_5396_8177.t157 a_n11317_n20927.t1 a_5396_n6451.t13 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X303 AVSS.t244 AVSS.t243 AVSS.t244 AVSS.t201 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X304 VOUT.t67 a_n11317_n20927.t1 a_5396_9163.t165 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X305 a_5396_9163.t72 a_5396_n6451.t97 AVDD.t1555 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X306 a_n13990_8177.t351 VN.t13 a_n13990_n5465.t99 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X307 AVSS.t242 AVSS.t241 AVSS.t242 AVSS.t133 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X308 AVDD.t1062 AVDD.t1061 AVDD.t1062 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X309 a_n13990_8177.t274 VP.t13 a_n13990_n6451.t128 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X310 a_n13990_n6451.t127 VP.t14 a_n13990_8177.t275 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X311 a_5396_9163.t164 a_n11317_n20927.t1 VOUT.t66 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X312 a_n13990_n6451.t126 VP.t15 a_n13990_8177.t276 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X313 AVDD.t1060 AVDD.t1059 AVDD.t1060 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X314 AVSS.t240 AVSS.t239 AVSS.t240 AVSS.t34 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X315 AVDD.t1058 AVDD.t1057 AVDD.t1058 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X316 a_n2101_n17634# a_n11317_n20927.t1 a_n2631_n17634# AVDD.t328 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X317 AVDD.t1056 AVDD.t1055 AVDD.t1056 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X318 a_n13990_8177.t288 VN.t14 a_n13990_n5465.t98 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X319 AVDD.t1556 a_5396_n6451.t98 a_5396_8177.t72 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X320 AVDD.t1054 AVDD.t1053 AVDD.t1054 AVDD.t153 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X321 a_n13990_8177.t289 VN.t15 a_n13990_n5465.t97 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X322 AVDD.t1690 IREF.t94 a_n13990_8177.t234 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X323 IREF.t33 IREF.t32 AVDD.t1599 AVDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X324 AVDD.t1052 AVDD.t1051 AVDD.t1052 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X325 AVDD.t1050 AVDD.t1049 AVDD.t1050 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X326 AVDD.t1048 AVDD.t1047 AVDD.t1048 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X327 AVDD.t1557 a_5396_n6451.t99 a_5396_9163.t71 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X328 AVDD.t1046 AVDD.t1045 AVDD.t1046 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X329 AVDD.t1044 AVDD.t1043 AVDD.t1044 AVDD.t638 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X330 AVSS.t238 AVSS.t237 AVSS.t238 AVSS.t43 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X331 AVDD.t1042 AVDD.t1041 AVDD.t1042 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X332 a_5396_9163.t70 a_5396_n6451.t100 AVDD.t1558 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X333 AVDD.t1040 AVDD.t1039 AVDD.t1040 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X334 a_n13990_n6451.t125 VP.t16 a_n13990_8177.t277 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X335 AVDD.t1559 a_5396_n6451.t101 a_5396_8177.t71 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X336 AVDD.t1038 AVDD.t1037 AVDD.t1038 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X337 AVDD.t1036 AVDD.t1035 AVDD.t1036 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X338 AVDD.t1034 AVDD.t1033 AVDD.t1034 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X339 IREF.t31 IREF.t30 AVDD.t1598 AVDD.t480 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X340 a_n13990_8177.t290 VN.t16 a_n13990_n5465.t96 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X341 AVDD.t1560 a_5396_n6451.t102 a_5396_8177.t70 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X342 AVDD.t1032 AVDD.t1031 AVDD.t1032 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X343 a_n13990_n5465.t95 VN.t17 a_n13990_8177.t291 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X344 AVDD.t1561 a_5396_n6451.t103 a_5396_9163.t69 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X345 a_5396_n6451.t12 a_n11317_n20927.t1 a_5396_8177.t156 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X346 VOUT.t65 a_n11317_n20927.t1 a_5396_9163.t103 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X347 a_5396_8177.t69 a_5396_n6451.t104 AVDD.t1562 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X348 AVDD.t1339 a_5396_n6451.t105 a_5396_8177.t68 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X349 a_5396_9163.t68 a_5396_n6451.t106 AVDD.t1340 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X350 AVSS.t236 AVSS.t234 AVSS.t236 AVSS.t235 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X351 AVDD.t1030 AVDD.t1029 AVDD.t1030 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X352 AVDD.t1563 IREF.t95 a_n13990_8177.t233 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X353 a_n13990_8177.t278 VP.t17 a_n13990_n6451.t124 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X354 a_n13990_n5465.t94 VN.t18 a_n13990_8177.t292 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X355 a_5396_n6451.t11 a_n11317_n20927.t1 a_5396_8177.t155 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X356 a_n13990_n6451.t123 VP.t18 a_n13990_8177.t307 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X357 AVDD.t1028 AVDD.t1027 AVDD.t1028 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X358 AVDD.t1026 AVDD.t1025 AVDD.t1026 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X359 a_5396_9163.t67 a_5396_n6451.t107 AVDD.t1341 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X360 AVDD.t1564 IREF.t96 a_n13990_8177.t232 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X361 a_n13990_n5465.t22 a_n11737_n14973.t41 AVSS.t335 AVSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X362 a_n13990_n5465.t129 a_n11737_n15980.t34 VOUT.t102 AVSS.t67 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X363 a_n13990_8177.t308 VP.t19 a_n13990_n6451.t122 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X364 a_n13990_n5465.t136 a_n11737_n15980.t35 VOUT.t101 AVSS.t64 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X365 a_n6139_n20820# a_n11737_n15980.t36 a_n6661_n21443# AVSS.t178 nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X366 AVDD.t1024 AVDD.t1023 AVDD.t1024 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X367 VOUT.t100 a_n11737_n15980.t37 a_n13990_n5465.t135 AVSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X368 a_n13990_8177.t309 VP.t20 a_n13990_n6451.t121 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X369 AVSS.t336 a_n11737_n14973.t42 a_n13990_n6451.t26 AVSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X370 AVDD.t1022 AVDD.t1021 AVDD.t1022 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X371 AVDD.t1565 IREF.t97 a_n11737_n14973.t24 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X372 AVDD.t1020 AVDD.t1019 AVDD.t1020 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X373 AVSS.t233 AVSS.t232 AVSS.t233 AVSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X374 a_n13990_8177.t310 VP.t21 a_n13990_n6451.t120 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X375 AVDD.t1018 AVDD.t1017 AVDD.t1018 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X376 a_n13990_n5465.t93 VN.t19 a_n13990_8177.t42 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X377 AVDD.t1016 AVDD.t1015 AVDD.t1016 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X378 AVDD.t1014 AVDD.t1013 AVDD.t1014 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X379 AVDD.t1012 AVDD.t1011 AVDD.t1012 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X380 a_n13990_8177.t311 VP.t22 a_n13990_n6451.t119 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X381 AVDD.t1010 AVDD.t1009 AVDD.t1010 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X382 AVDD.t1566 IREF.t98 a_n13990_8177.t231 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X383 AVDD.t1342 a_5396_n6451.t108 a_5396_9163.t66 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X384 AVDD.t1008 AVDD.t1007 AVDD.t1008 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X385 AVDD.t1597 IREF.t28 IREF.t29 AVDD.t282 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X386 a_n13990_8177.t43 VN.t20 a_n13990_n5465.t92 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X387 AVDD.t1343 a_5396_n6451.t109 a_5396_8177.t67 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X388 AVDD.t1567 IREF.t99 a_n13990_8177.t230 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X389 AVDD.t1006 AVDD.t1005 AVDD.t1006 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X390 AVDD.t1004 AVDD.t1003 AVDD.t1004 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X391 AVDD.t1568 IREF.t100 a_n11737_n15980.t17 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X392 AVSS.t337 a_n11737_n14973.t43 a_n13990_n6451.t27 AVSS.t82 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X393 a_n965_n16909# a_n11317_n20927.t1 a_n1533_n16909# AVDD.t264 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X394 a_5396_9163.t102 a_n11317_n20927.t1 VOUT.t64 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X395 AVDD.t1002 AVDD.t1001 AVDD.t1002 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X396 a_5396_8177.t154 a_n11317_n20927.t1 a_5396_n6451.t10 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X397 AVDD.t1000 AVDD.t999 AVDD.t1000 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X398 a_n13990_8177.t44 VN.t21 a_n13990_n5465.t91 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X399 AVDD.t998 AVDD.t997 AVDD.t998 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X400 AVDD.t996 AVDD.t995 AVDD.t996 AVDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X401 AVDD.t1344 a_5396_n6451.t110 a_5396_9163.t65 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X402 a_n13990_n6451.t118 VP.t23 a_n13990_8177.t93 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X403 AVDD.t994 AVDD.t993 AVDD.t994 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X404 AVSS.t231 AVSS.t230 AVSS.t231 AVSS.t25 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X405 AVDD.t1345 a_5396_n6451.t111 a_5396_8177.t66 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X406 a_5396_8177.t153 a_n11317_n20927.t1 a_5396_n6451.t9 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X407 a_5396_8177.t65 a_5396_n6451.t112 AVDD.t1346 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X408 AVSS.t229 AVSS.t228 AVSS.t229 AVSS.t28 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X409 a_5396_9163.t93 a_n11317_n20927.t1 VOUT.t63 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X410 a_5396_8177.t152 a_n11317_n20927.t1 a_5396_n6451.t8 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X411 AVDD.t1569 IREF.t101 a_n13990_8177.t229 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X412 AVDD.t992 AVDD.t991 AVDD.t992 AVDD.t2 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X413 a_5396_n6451.t7 a_n11317_n20927.t1 a_5396_8177.t151 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X414 AVDD.t990 AVDD.t989 AVDD.t990 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X415 a_5396_n6451.t6 a_n11317_n20927.t1 a_5396_8177.t150 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X416 AVDD.t988 AVDD.t987 AVDD.t988 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X417 AVDD.t1570 IREF.t102 a_n13990_8177.t228 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X418 a_5396_8177.t149 a_n11317_n20927.t1 a_5396_n6451.t5 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X419 AVDD.t986 AVDD.t985 AVDD.t986 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X420 AVSS.t363 a_n11737_n14973.t6 a_n11737_n14973.t7 AVSS.t138 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X421 a_n13990_8177.t45 VN.t22 a_n13990_n5465.t90 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X422 AVSS.t227 AVSS.t226 AVSS.t227 AVSS.t175 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X423 a_5396_n6451.t53 a_n11317_n20927.t1 a_5396_8177.t148 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X424 AVDD.t984 AVDD.t983 AVDD.t984 AVDD.t181 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X425 AVSS.t225 AVSS.t224 AVSS.t225 AVSS.t172 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X426 AVDD.t982 AVDD.t981 AVDD.t982 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X427 a_n13990_8177.t227 IREF.t103 AVDD.t1571 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X428 a_n13990_8177.t226 IREF.t104 AVDD.t1572 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X429 AVDD.t980 AVDD.t979 AVDD.t980 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X430 AVSS.t348 a_n11737_n14973.t44 a_n13990_n5465.t118 AVSS.t114 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X431 VOUT.t62 a_n11317_n20927.t1 a_5396_9163.t92 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X432 a_5396_9163.t141 a_n11317_n20927.t1 VOUT.t61 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X433 AVDD.t978 AVDD.t977 AVDD.t978 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X434 a_n13990_n6451.t117 VP.t24 a_n13990_8177.t94 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X435 a_5396_8177.t147 a_n11317_n20927.t1 a_5396_n6451.t35 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X436 AVDD.t976 AVDD.t975 AVDD.t976 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X437 AVDD.t974 AVDD.t973 AVDD.t974 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X438 a_5396_8177.t64 a_5396_n6451.t113 AVDD.t1347 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X439 a_5396_8177.t63 a_5396_n6451.t114 AVDD.t1348 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X440 AVDD.t972 AVDD.t971 AVDD.t972 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X441 a_n13990_8177.t46 VN.t23 a_n13990_n5465.t89 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X442 a_n13990_8177.t225 IREF.t105 AVDD.t1573 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X443 AVDD.t970 AVDD.t969 AVDD.t970 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X444 AVSS.t223 AVSS.t221 AVSS.t223 AVSS.t222 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X445 AVDD.t968 AVDD.t967 AVDD.t968 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X446 a_n11737_n14973.t23 IREF.t106 AVDD.t1574 AVDD.t39 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X447 AVDD.t966 AVDD.t965 AVDD.t966 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X448 AVSS.t349 a_n11737_n14973.t45 a_n13990_n5465.t119 AVSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X449 AVSS.t350 a_n11737_n14973.t46 a_n13990_n6451.t30 AVSS.t19 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X450 AVSS.t351 a_n11737_n14973.t47 a_n13990_n5465.t120 AVSS.t16 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X451 AVDD.t964 AVDD.t963 AVDD.t964 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X452 AVDD.t962 AVDD.t961 AVDD.t962 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X453 a_5396_n6451.t64 a_n11737_n15980.t38 a_n13990_n6451.t42 AVSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X454 AVSS.t317 a_n11737_n14973.t48 a_n11317_n20927.t1 AVSS.t133 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X455 AVDD.t960 AVDD.t959 AVDD.t960 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X456 a_5396_n6451.t65 a_n11737_n15980.t39 a_n13990_n6451.t41 AVSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X457 AVDD.t958 AVDD.t957 AVDD.t958 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X458 AVDD.t956 AVDD.t955 AVDD.t956 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X459 AVSS.t220 AVSS.t219 AVSS.t220 AVSS.t88 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X460 AVSS.t218 AVSS.t217 AVSS.t218 AVSS.t85 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X461 a_n11737_n14973.t22 IREF.t107 AVDD.t1575 AVDD.t480 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X462 a_n13990_n6451.t116 VP.t25 a_n13990_8177.t95 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X463 a_n13990_8177.t96 VP.t26 a_n13990_n6451.t115 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X464 a_n13990_8177.t97 VP.t27 a_n13990_n6451.t114 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X465 AVDD.t954 AVDD.t953 AVDD.t954 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X466 a_n13990_n6451.t113 VP.t28 a_n13990_8177.t298 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X467 AVDD.t952 AVDD.t951 AVDD.t952 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X468 VOUT.t60 a_n11317_n20927.t1 a_5396_9163.t140 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X469 AVDD.t950 AVDD.t949 AVDD.t950 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X470 a_5396_n6451.t52 a_n11317_n20927.t1 a_5396_8177.t146 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X471 a_n13990_n6451.t112 VP.t29 a_n13990_8177.t299 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X472 a_5396_8177.t62 a_5396_n6451.t115 AVDD.t1349 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X473 a_5396_8177.t61 a_5396_n6451.t116 AVDD.t1350 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X474 a_n13990_n5465.t88 VN.t24 a_n13990_8177.t37 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X475 AVDD.t1351 a_5396_n6451.t117 a_5396_9163.t64 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X476 AVDD.t948 AVDD.t947 AVDD.t948 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X477 a_n11737_n15980.t16 IREF.t108 AVDD.t1576 AVDD.t480 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X478 AVDD.t1577 IREF.t109 a_n13990_8177.t224 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X479 a_5396_9163.t63 a_5396_n6451.t118 AVDD.t1352 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X480 AVDD.t946 AVDD.t945 AVDD.t946 AVDD.t131 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X481 VOUT.t59 a_n11317_n20927.t1 a_5396_9163.t129 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X482 AVDD.t944 AVDD.t943 AVDD.t944 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X483 AVDD.t942 AVDD.t941 AVDD.t942 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X484 a_n13990_8177.t223 IREF.t110 AVDD.t1578 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X485 a_5396_n6451.t52 a_n11317_n20927.t1 a_5396_8177.t145 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X486 AVDD.t1353 a_5396_n6451.t119 a_5396_9163.t62 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X487 AVDD.t940 AVDD.t939 AVDD.t940 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X488 AVDD.t938 AVDD.t937 AVDD.t938 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X489 AVDD.t936 AVDD.t935 AVDD.t936 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X490 AVDD.t934 AVDD.t933 AVDD.t934 AVDD.t178 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X491 AVSS.t216 AVSS.t215 AVSS.t216 AVSS.t49 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X492 a_n13990_8177.t38 VN.t25 a_n13990_n5465.t87 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X493 a_n13990_n6451.t111 VP.t30 a_n13990_8177.t300 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X494 AVSS.t318 a_n11737_n14973.t49 a_n13990_n5465.t13 AVSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X495 a_n13990_8177.t222 IREF.t111 AVDD.t1579 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X496 AVDD.t932 AVDD.t931 AVDD.t932 AVDD.t13 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X497 AVDD.t1657 IREF.t112 a_n13990_8177.t221 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X498 AVDD.t930 AVDD.t929 AVDD.t930 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X499 AVDD.t1658 IREF.t113 a_n13990_8177.t220 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X500 a_5396_8177.t60 a_5396_n6451.t120 AVDD.t1354 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X501 a_n13990_8177.t219 IREF.t114 AVDD.t1659 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X502 AVSS.t214 AVSS.t213 AVSS.t214 AVSS.t79 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X503 AVSS.t212 AVSS.t211 AVSS.t212 AVSS.t31 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X504 AVDD.t1660 IREF.t115 a_n13990_8177.t218 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X505 a_n13990_8177.t39 VN.t26 a_n13990_n5465.t86 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X506 AVSS.t210 AVSS.t209 AVSS.t210 AVSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X507 a_n13990_n6451.t110 VP.t31 a_n13990_8177.t301 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X508 AVDD.t928 AVDD.t927 AVDD.t928 AVDD.t156 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X509 AVDD.t926 AVDD.t925 AVDD.t926 AVDD.t27 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X510 AVDD.t924 AVDD.t923 AVDD.t924 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X511 AVDD.t922 AVDD.t921 AVDD.t922 AVDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X512 a_n13990_8177.t40 VN.t27 a_n13990_n5465.t85 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X513 a_5396_8177.t144 a_n11317_n20927.t1 a_5396_n6451.t44 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X514 AVDD.t1355 a_5396_n6451.t121 a_5396_8177.t59 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X515 AVDD.t920 AVDD.t919 AVDD.t920 AVDD.t373 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X516 AVSS.t208 AVSS.t207 AVSS.t208 AVSS.t158 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X517 AVSS.t206 AVSS.t205 AVSS.t206 AVSS.t155 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X518 AVSS.t204 AVSS.t203 AVSS.t204 AVSS.t46 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X519 AVDD.t918 AVDD.t917 AVDD.t918 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X520 a_5396_9163.t61 a_5396_n6451.t122 AVDD.t1356 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X521 AVDD.t916 AVDD.t915 AVDD.t916 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X522 AVDD.t914 AVDD.t913 AVDD.t914 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X523 a_n13990_8177.t41 VN.t28 a_n13990_n5465.t84 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X524 a_n13990_n6451.t109 VP.t32 a_n13990_8177.t302 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X525 a_5396_n6451.t47 a_n11317_n20927.t1 a_5396_8177.t143 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X526 AVDD.t912 AVDD.t911 AVDD.t912 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X527 AVDD.t910 AVDD.t909 AVDD.t910 AVDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X528 AVDD.t908 AVDD.t907 AVDD.t908 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X529 a_n13990_8177.t32 VN.t29 a_n13990_n5465.t83 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X530 a_5396_n6451.t62 a_n11317_n20927.t4 a_5396_8177.t175 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X531 a_n13990_8177.t217 IREF.t116 AVDD.t1661 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X532 AVDD.t906 AVDD.t905 AVDD.t906 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X533 AVDD.t904 AVDD.t903 AVDD.t904 AVDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X534 AVSS.t202 AVSS.t200 AVSS.t202 AVSS.t201 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X535 a_5396_8177.t58 a_5396_n6451.t123 AVDD.t1357 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X536 AVSS.t199 AVSS.t198 AVSS.t199 AVSS.t67 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X537 a_5396_9163.t60 a_5396_n6451.t124 AVDD.t1358 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X538 AVSS.t197 AVSS.t196 AVSS.t197 AVSS.t64 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X539 AVDD.t902 AVDD.t901 AVDD.t902 AVDD.t480 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X540 a_n13990_n5465.t82 VN.t30 a_n13990_8177.t33 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X541 IREF.t27 IREF.t26 AVDD.t1699 AVDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X542 a_n13990_8177.t216 IREF.t117 AVDD.t1662 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X543 AVDD.t900 AVDD.t899 AVDD.t900 AVDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X544 a_5396_n6451.t47 a_n11317_n20927.t1 a_5396_8177.t142 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X545 AVSS.t319 a_n11737_n14973.t50 a_n13990_n5465.t14 AVSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X546 a_5396_9163.t128 a_n11317_n20927.t1 VOUT.t58 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X547 a_5396_9163.t117 a_n11317_n20927.t1 VOUT.t57 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X548 AVDD.t898 AVDD.t897 AVDD.t898 AVDD.t13 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X549 a_n13990_n5465.t122 a_n11737_n15980.t40 VOUT.t99 AVSS.t37 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X550 VOUT.t56 a_n11317_n20927.t1 a_5396_9163.t116 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X551 a_5396_9163.t131 a_n11317_n20927.t1 VOUT.t55 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X552 AVDD.t1359 a_5396_n6451.t125 a_5396_8177.t57 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X553 AVDD.t896 AVDD.t895 AVDD.t896 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X554 AVSS.t195 AVSS.t194 AVSS.t195 AVSS.t43 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X555 a_n13990_n5465.t81 VN.t31 a_n13990_8177.t34 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X556 AVDD.t894 AVDD.t893 AVDD.t894 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X557 AVDD.t892 AVDD.t891 AVDD.t892 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X558 AVDD.t1360 a_5396_n6451.t126 a_5396_9163.t59 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X559 AVDD.t890 AVDD.t889 AVDD.t890 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X560 AVDD.t1361 a_5396_n6451.t127 a_5396_9163.t58 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X561 AVDD.t1362 a_5396_n6451.t128 a_5396_8177.t56 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X562 a_5396_8177.t141 a_n11317_n20927.t1 a_5396_n6451.t51 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X563 a_5396_9163.t130 a_n11317_n20927.t1 VOUT.t54 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X564 AVDD.t1663 IREF.t118 a_n11737_n14973.t21 AVDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X565 AVDD.t888 AVDD.t887 AVDD.t888 AVDD.t373 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X566 VOUT.t53 a_n11317_n20927.t1 a_5396_9163.t111 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X567 a_5396_9163.t110 a_n11317_n20927.t1 VOUT.t52 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X568 AVDD.t886 AVDD.t885 AVDD.t886 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X569 AVDD.t1664 IREF.t119 a_n13990_8177.t215 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X570 AVDD.t884 AVDD.t883 AVDD.t884 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X571 AVSS.t193 AVSS.t192 AVSS.t193 AVSS.t34 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X572 a_n13990_8177.t337 VP.t33 a_n13990_n6451.t108 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X573 a_5396_9163.t161 a_n11317_n20927.t1 VOUT.t51 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X574 a_5396_n6451.t50 a_n11317_n20927.t1 a_5396_8177.t140 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X575 AVDD.t882 AVDD.t881 AVDD.t882 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X576 AVDD.t880 AVDD.t879 AVDD.t880 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X577 AVDD.t878 AVDD.t877 AVDD.t878 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X578 a_n13990_8177.t214 IREF.t120 AVDD.t1665 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X579 a_n13990_n6451.t20 a_n11737_n14973.t51 AVSS.t320 AVSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X580 a_n13990_n6451.t9 a_n11737_n14973.t52 AVSS.t295 AVSS.t16 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X581 AVSS.t296 a_n11737_n14973.t53 a_n13990_n5465.t3 AVSS.t19 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X582 VOUT.t98 a_n11737_n15980.t41 a_n13990_n5465.t121 AVSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X583 a_5396_8177.t55 a_5396_n6451.t129 AVDD.t1363 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X584 VOUT.t97 a_n11737_n15980.t42 a_n13990_n5465.t132 AVSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X585 AVDD.t876 AVDD.t874 AVDD.t876 AVDD.t875 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X586 a_n13990_8177.t35 VN.t32 a_n13990_n5465.t80 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X587 a_5396_9163.t160 a_n11317_n20927.t1 VOUT.t50 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X588 AVDD.t873 AVDD.t872 AVDD.t873 AVDD.t178 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X589 a_n13990_n5465.t79 VN.t33 a_n13990_8177.t36 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X590 AVSS.t191 AVSS.t190 AVSS.t191 AVSS.t144 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X591 a_5396_9163.t57 a_5396_n6451.t130 AVDD.t1364 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X592 AVSS.t189 AVSS.t188 AVSS.t189 AVSS.t141 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X593 AVDD.t871 AVDD.t870 AVDD.t871 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X594 AVDD.t869 AVDD.t868 AVDD.t869 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X595 AVDD.t1666 IREF.t121 a_n11737_n14973.t20 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X596 AVDD.t867 AVDD.t866 AVDD.t867 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X597 AVDD.t865 AVDD.t864 AVDD.t865 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X598 AVDD.t863 AVDD.t862 AVDD.t863 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X599 AVDD.t861 AVDD.t860 AVDD.t861 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X600 AVDD.t1365 a_5396_n6451.t131 a_5396_8177.t54 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X601 a_n13990_8177.t213 IREF.t122 AVDD.t1667 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X602 AVSS.t187 AVSS.t186 AVSS.t187 AVSS.t178 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X603 a_n13990_8177.t212 IREF.t123 AVDD.t1668 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X604 AVDD.t859 AVDD.t858 AVDD.t859 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X605 AVDD.t857 AVDD.t856 AVDD.t857 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X606 AVDD.t855 AVDD.t854 AVDD.t855 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X607 a_n13990_n5465.t78 VN.t34 a_n13990_8177.t27 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X608 AVDD.t1698 IREF.t24 IREF.t25 AVDD.t282 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X609 AVDD.t853 AVDD.t852 AVDD.t853 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X610 AVDD.t851 AVDD.t850 AVDD.t851 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X611 AVDD.t849 AVDD.t848 AVDD.t849 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X612 a_5396_9163.t56 a_5396_n6451.t132 AVDD.t1366 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X613 a_n13990_n6451.t10 a_n11737_n14973.t54 AVSS.t297 AVSS.t235 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X614 a_n13990_8177.t211 IREF.t124 AVDD.t1669 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X615 a_5396_9163.t55 a_5396_n6451.t133 AVDD.t1367 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X616 AVSS.t298 a_n11737_n14973.t55 a_n13990_n5465.t4 AVSS.t82 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X617 AVDD.t847 AVDD.t846 AVDD.t847 AVDD.t193 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X618 AVDD.t845 AVDD.t844 AVDD.t845 AVDD.t178 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X619 AVDD.t843 AVDD.t842 AVDD.t843 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X620 AVDD.t841 AVDD.t840 AVDD.t841 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X621 AVDD.t839 AVDD.t838 AVDD.t839 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X622 a_5396_n6451.t2 a_n11737_n15980.t43 a_n13990_n6451.t40 AVSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X623 AVDD.t1368 a_5396_n6451.t134 a_5396_8177.t53 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X624 a_n13990_8177.t210 IREF.t125 AVDD.t1670 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X625 AVDD.t837 AVDD.t836 AVDD.t837 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X626 AVDD.t835 AVDD.t834 AVDD.t835 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X627 a_5396_9163.t113 a_n11317_n20927.t1 VOUT.t49 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X628 AVDD.t833 AVDD.t832 AVDD.t833 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X629 AVDD.t831 AVDD.t830 AVDD.t831 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X630 AVDD.t829 AVDD.t828 AVDD.t829 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X631 a_n13990_8177.t209 IREF.t126 AVDD.t1671 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X632 AVDD.t827 AVDD.t826 AVDD.t827 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X633 a_n13990_8177.t208 IREF.t127 AVDD.t1672 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X634 AVSS.t185 AVSS.t184 AVSS.t185 AVSS.t25 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X635 AVDD.t825 AVDD.t824 AVDD.t825 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X636 a_n13990_8177.t207 IREF.t128 AVDD.t1673 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X637 AVDD.t823 AVDD.t822 AVDD.t823 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X638 AVDD.t1286 IREF.t129 a_n13990_8177.t206 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X639 a_n11737_n15980.t15 IREF.t130 AVDD.t1287 AVDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X640 AVDD.t821 AVDD.t820 AVDD.t821 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X641 AVDD.t1369 a_5396_n6451.t135 a_5396_9163.t54 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X642 a_n13990_8177.t205 IREF.t131 AVDD.t1288 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X643 a_n13990_8177.t338 VP.t34 a_n13990_n6451.t107 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X644 AVDD.t819 AVDD.t818 AVDD.t819 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X645 AVDD.t817 AVDD.t816 AVDD.t817 AVDD.t181 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X646 AVSS.t183 AVSS.t182 AVSS.t183 AVSS.t79 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X647 AVDD.t815 AVDD.t814 AVDD.t815 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X648 IREF.t23 IREF.t22 AVDD.t1697 AVDD.t39 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X649 a_5396_8177.t52 a_5396_n6451.t136 AVDD.t1370 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X650 AVDD.t1289 IREF.t132 a_n13990_8177.t204 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X651 AVDD.t1371 a_5396_n6451.t137 a_5396_9163.t53 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X652 AVSS.t181 AVSS.t180 AVSS.t181 AVSS.t95 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X653 AVDD.t813 AVDD.t812 AVDD.t813 AVDD.t153 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X654 AVDD.t811 AVDD.t809 AVDD.t811 AVDD.t810 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X655 AVDD.t808 AVDD.t807 AVDD.t808 AVDD.t2 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X656 AVSS.t179 AVSS.t177 AVSS.t179 AVSS.t178 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X657 a_n11737_n14973.t19 IREF.t133 AVDD.t1290 AVDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X658 AVDD.t806 AVDD.t805 AVDD.t806 AVDD.t13 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X659 AVSS.t176 AVSS.t174 AVSS.t176 AVSS.t175 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X660 AVSS.t173 AVSS.t171 AVSS.t173 AVSS.t172 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X661 VOUT.t48 a_n11317_n20927.t1 a_5396_9163.t112 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X662 AVDD.t804 AVDD.t803 AVDD.t804 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X663 a_n965_n15598# a_n11317_n20927.t1 a_n1533_n15598# AVDD.t264 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X664 AVDD.t802 AVDD.t801 AVDD.t802 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X665 AVDD.t800 AVDD.t799 AVDD.t800 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X666 a_5396_8177.t51 a_5396_n6451.t138 AVDD.t1372 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X667 a_5396_8177.t50 a_5396_n6451.t139 AVDD.t1373 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X668 a_n13990_n6451.t106 VP.t35 a_n13990_8177.t339 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X669 AVDD.t798 AVDD.t797 AVDD.t798 AVDD.t373 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X670 a_n11737_n15980.t14 IREF.t134 AVDD.t1291 AVDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X671 AVDD.t796 AVDD.t795 AVDD.t796 AVDD.t156 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X672 a_n13990_8177.t203 IREF.t135 AVDD.t1292 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X673 a_n13990_8177.t202 IREF.t136 AVDD.t1293 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X674 AVDD.t794 AVDD.t793 AVDD.t794 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X675 AVDD.t1294 IREF.t137 a_n13990_8177.t201 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X676 AVDD.t1304 a_5396_n6451.t140 a_5396_9163.t52 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X677 AVDD.t792 AVDD.t791 AVDD.t792 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X678 AVDD.t790 AVDD.t789 AVDD.t790 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X679 AVDD.t788 AVDD.t787 AVDD.t788 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X680 a_5396_8177.t49 a_5396_n6451.t141 AVDD.t1305 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X681 a_5396_9163.t51 a_5396_n6451.t142 AVDD.t1306 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X682 AVDD.t1295 IREF.t138 a_n13990_8177.t200 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X683 AVDD.t786 AVDD.t785 AVDD.t786 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X684 a_5396_8177.t139 a_n11317_n20927.t1 a_5396_n6451.t40 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X685 VOUT.t47 a_n11317_n20927.t1 a_5396_9163.t107 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X686 a_n13990_8177.t28 VN.t35 a_n13990_n5465.t77 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X687 AVSS.t170 AVSS.t169 AVSS.t170 AVSS.t74 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X688 AVDD.t784 AVDD.t783 AVDD.t784 AVDD.t131 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X689 a_n13990_n6451.t52 a_n11737_n14973.t56 AVSS.t358 AVSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X690 AVDD.t782 AVDD.t781 AVDD.t782 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X691 AVDD.t1307 a_5396_n6451.t143 a_5396_9163.t50 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X692 a_n13990_n6451.t105 VP.t36 a_n13990_8177.t340 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X693 a_n13990_8177.t199 IREF.t139 AVDD.t1296 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X694 a_n13990_8177.t198 IREF.t140 AVDD.t1297 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X695 AVDD.t780 AVDD.t779 AVDD.t780 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X696 AVDD.t778 AVDD.t777 AVDD.t778 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X697 a_5396_8177.t138 a_n11317_n20927.t1 a_5396_n6451.t39 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X698 a_n13990_n6451.t104 VP.t37 a_n13990_8177.t341 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X699 AVDD.t776 AVDD.t775 AVDD.t776 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X700 a_n13990_n5465.t140 a_n11737_n14973.t57 AVSS.t359 AVSS.t222 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X701 VOUT.t46 a_n11317_n20927.t1 a_5396_9163.t106 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X702 AVDD.t774 AVDD.t773 AVDD.t774 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X703 AVDD.t772 AVDD.t771 AVDD.t772 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X704 AVDD.t1298 IREF.t141 a_n11737_n15980.t13 AVDD.t810 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X705 a_n13990_8177.t197 IREF.t142 AVDD.t1299 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X706 AVDD.t1300 IREF.t143 a_n13990_8177.t196 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X707 AVDD.t1301 IREF.t144 a_n13990_8177.t195 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X708 a_5396_n6451.t38 a_n11317_n20927.t1 a_5396_8177.t137 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X709 AVDD.t770 AVDD.t769 AVDD.t770 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X710 AVDD.t768 AVDD.t767 AVDD.t768 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X711 AVDD.t766 AVDD.t765 AVDD.t766 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X712 AVDD.t764 AVDD.t763 AVDD.t764 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X713 a_5396_n6451.t37 a_n11317_n20927.t1 a_5396_8177.t136 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X714 a_n13990_n6451.t103 VP.t38 a_n13990_8177.t293 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X715 a_n965_n16909# a_n11317_n20927.t1 a_n1533_n16323# AVDD.t264 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X716 AVSS.t168 AVSS.t167 AVSS.t168 AVSS.t49 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X717 AVDD.t762 AVDD.t761 AVDD.t762 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X718 AVDD.t1302 IREF.t145 a_n11737_n14973.t18 AVDD.t282 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X719 a_5396_9163.t169 a_n11317_n20927.t1 VOUT.t45 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X720 AVDD.t1303 IREF.t146 a_n13990_8177.t194 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X721 AVDD.t760 AVDD.t759 AVDD.t760 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X722 AVDD.t758 AVDD.t757 AVDD.t758 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X723 a_5396_8177.t48 a_5396_n6451.t144 AVDD.t1308 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X724 AVDD.t756 AVDD.t755 AVDD.t756 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X725 AVDD.t754 AVDD.t753 AVDD.t754 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X726 AVDD.t752 AVDD.t751 AVDD.t752 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X727 AVDD.t750 AVDD.t749 AVDD.t750 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X728 AVSS.t360 a_n11737_n14973.t58 a_n13990_n5465.t141 AVSS.t235 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X729 AVSS.t166 AVSS.t165 AVSS.t166 AVSS.t37 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X730 a_n13990_n6451.t102 VP.t39 a_n13990_8177.t294 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X731 a_n11737_n14973.t5 a_n11737_n14973.t4 AVSS.t362 AVSS.t31 nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X732 AVSS.t164 AVSS.t162 AVSS.t164 AVSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X733 AVDD.t748 AVDD.t747 AVDD.t748 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X734 AVDD.t746 AVDD.t745 AVDD.t746 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X735 a_5396_8177.t47 a_5396_n6451.t145 AVDD.t1309 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X736 AVDD.t744 AVDD.t743 AVDD.t744 AVDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X737 AVDD.t1310 a_5396_n6451.t146 a_5396_9163.t49 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X738 a_n13990_8177.t193 IREF.t147 AVDD.t1459 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X739 a_n13990_8177.t192 IREF.t148 AVDD.t1460 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X740 AVDD.t742 AVDD.t741 AVDD.t742 AVDD.t394 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X741 AVDD.t740 AVDD.t739 AVDD.t740 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X742 AVDD.t738 AVDD.t737 AVDD.t738 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X743 AVSS.t161 AVSS.t160 AVSS.t161 AVSS.t55 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X744 AVSS.t159 AVSS.t157 AVSS.t159 AVSS.t158 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X745 AVDD.t736 AVDD.t735 AVDD.t736 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X746 AVDD.t734 AVDD.t733 AVDD.t734 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X747 AVSS.t156 AVSS.t154 AVSS.t156 AVSS.t155 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X748 a_5396_n6451.t36 a_n11317_n20927.t1 a_5396_8177.t135 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X749 AVDD.t1461 IREF.t149 a_n11737_n15980.t12 AVDD.t282 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X750 a_n13990_8177.t191 IREF.t150 AVDD.t1462 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X751 AVSS.t153 AVSS.t152 AVSS.t153 AVSS.t13 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X752 a_n13990_n5465.t76 VN.t36 a_n13990_8177.t29 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X753 a_5396_8177.t46 a_5396_n6451.t147 AVDD.t1311 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X754 AVSS.t151 AVSS.t150 AVSS.t151 AVSS.t10 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X755 a_5396_n6451.t10 a_n11317_n20927.t1 a_5396_8177.t134 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X756 AVSS.t149 AVSS.t148 AVSS.t149 AVSS.t34 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X757 AVDD.t732 AVDD.t731 AVDD.t732 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X758 AVSS.t333 a_n11737_n15980.t44 a_n6139_n21443# AVSS.t98 nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X759 AVDD.t730 AVDD.t729 AVDD.t730 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X760 AVDD.t728 AVDD.t727 AVDD.t728 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X761 AVSS.t361 a_n11737_n14973.t59 a_n13990_n6451.t53 AVSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X762 a_n13990_n5465.t131 a_n11737_n15980.t45 VOUT.t96 AVSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X763 AVDD.t726 AVDD.t725 AVDD.t726 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X764 AVDD.t724 AVDD.t723 AVDD.t724 AVDD.t181 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X765 AVDD.t722 AVDD.t721 AVDD.t722 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X766 AVDD.t720 AVDD.t719 AVDD.t720 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X767 AVDD.t718 AVDD.t716 AVDD.t718 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X768 a_5396_n6451.t9 a_n11317_n20927.t1 a_5396_8177.t133 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X769 AVDD.t715 AVDD.t714 AVDD.t715 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X770 AVDD.t713 AVDD.t712 AVDD.t713 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X771 a_n13990_8177.t190 IREF.t151 AVDD.t1463 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X772 AVDD.t711 AVDD.t710 AVDD.t711 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X773 a_n13990_8177.t189 IREF.t152 AVDD.t1464 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X774 a_5396_9163.t48 a_5396_n6451.t148 AVDD.t1312 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X775 a_n13990_8177.t295 VP.t40 a_n13990_n6451.t101 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X776 AVDD.t709 AVDD.t708 AVDD.t709 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X777 AVDD.t707 AVDD.t706 AVDD.t707 AVDD.t181 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X778 AVDD.t705 AVDD.t704 AVDD.t705 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X779 AVDD.t1696 IREF.t20 IREF.t21 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X780 a_5396_9163.t47 a_5396_n6451.t149 AVDD.t1313 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X781 AVDD.t1465 IREF.t153 a_n13990_8177.t188 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X782 AVDD.t703 AVDD.t702 AVDD.t703 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X783 a_5396_8177.t45 a_5396_n6451.t150 AVDD.t1314 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X784 a_n13990_n6451.t22 a_n11737_n14973.t60 AVSS.t329 AVSS.t201 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X785 AVDD.t701 AVDD.t700 AVDD.t701 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X786 AVDD.t699 AVDD.t698 AVDD.t699 AVDD.t193 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X787 AVDD.t1466 IREF.t154 a_n13990_8177.t187 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X788 AVDD.t697 AVDD.t696 AVDD.t697 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X789 AVDD.t695 AVDD.t694 AVDD.t695 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X790 AVDD.t693 AVDD.t692 AVDD.t693 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X791 a_5396_8177.t132 a_n11317_n20927.t1 a_5396_n6451.t12 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X792 a_n11737_n14973.t3 a_n11737_n14973.t2 AVSS.t353 AVSS.t95 nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X793 AVDD.t691 AVDD.t690 AVDD.t691 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X794 AVDD.t689 AVDD.t688 AVDD.t689 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X795 a_n13990_n6451.t100 VP.t41 a_n13990_8177.t296 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X796 a_n13990_n5465.t75 VN.t37 a_n13990_8177.t30 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X797 AVDD.t687 AVDD.t686 AVDD.t687 AVDD.t282 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X798 AVDD.t685 AVDD.t684 AVDD.t685 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X799 AVDD.t683 AVDD.t682 AVDD.t683 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X800 AVDD.t1315 a_5396_n6451.t151 a_5396_8177.t44 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X801 VOUT.t44 a_n11317_n20927.t1 a_5396_9163.t168 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X802 AVDD.t1316 a_5396_n6451.t152 a_5396_9163.t46 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X803 a_5396_8177.t43 a_5396_n6451.t153 AVDD.t1317 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X804 AVSS.t147 AVSS.t146 AVSS.t147 AVSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X805 AVDD.t681 AVDD.t680 AVDD.t681 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X806 a_n13990_8177.t186 IREF.t155 AVDD.t1467 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X807 a_5396_9163.t139 a_n11317_n20927.t1 VOUT.t43 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X808 a_n13990_n6451.t99 VP.t42 a_n13990_8177.t297 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X809 a_n13990_n5465.t74 VN.t38 a_n13990_8177.t31 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X810 AVDD.t679 AVDD.t678 AVDD.t679 AVDD.t131 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X811 AVDD.t677 AVDD.t676 AVDD.t677 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X812 AVSS.t145 AVSS.t143 AVSS.t145 AVSS.t144 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X813 AVSS.t142 AVSS.t140 AVSS.t142 AVSS.t141 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X814 AVDD.t675 AVDD.t674 AVDD.t675 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X815 AVDD.t673 AVDD.t672 AVDD.t673 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X816 AVDD.t671 AVDD.t670 AVDD.t671 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X817 AVDD.t669 AVDD.t668 AVDD.t669 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X818 AVDD.t667 AVDD.t666 AVDD.t667 AVDD.t328 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X819 AVDD.t1468 IREF.t156 a_n13990_8177.t185 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X820 AVDD.t1318 a_5396_n6451.t154 a_5396_9163.t45 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X821 AVDD.t1469 IREF.t157 a_n13990_8177.t184 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X822 AVDD.t1319 a_5396_n6451.t155 a_5396_8177.t42 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X823 AVDD.t665 AVDD.t664 AVDD.t665 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X824 AVDD.t1470 IREF.t158 a_n13990_8177.t183 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X825 AVDD.t663 AVDD.t662 AVDD.t663 AVDD.t153 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X826 AVDD.t1320 a_5396_n6451.t156 a_5396_8177.t41 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X827 a_n11737_n14973.t17 IREF.t159 AVDD.t1471 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X828 a_5396_9163.t44 a_5396_n6451.t157 AVDD.t1321 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X829 AVSS.t330 a_n11737_n14973.t61 a_n13990_n6451.t23 AVSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X830 AVDD.t661 AVDD.t660 AVDD.t661 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X831 AVSS.t331 a_n11737_n14973.t62 a_n13990_n6451.t24 AVSS.t222 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X832 a_5396_n6451.t35 a_n11317_n20927.t1 a_5396_8177.t131 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X833 a_5396_9163.t138 a_n11317_n20927.t1 VOUT.t42 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X834 a_5396_n6451.t34 a_n11317_n20927.t1 a_5396_8177.t130 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X835 a_n13990_n6451.t98 VP.t43 a_n13990_8177.t283 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X836 AVDD.t659 AVDD.t658 AVDD.t659 AVDD.t131 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X837 AVDD.t1322 a_5396_n6451.t158 a_5396_9163.t43 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X838 AVDD.t1379 a_n11317_n20927.t1 a_n1533_n17634# AVDD.t264 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X839 AVDD.t657 AVDD.t656 AVDD.t657 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X840 AVDD.t655 AVDD.t654 AVDD.t655 AVDD.t181 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X841 VOUT.t41 a_n11317_n20927.t1 a_5396_9163.t89 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X842 AVDD.t653 AVDD.t652 AVDD.t653 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X843 AVDD.t651 AVDD.t650 AVDD.t651 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X844 a_n13990_n5465.t73 VN.t39 a_n13990_8177.t22 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X845 a_n13990_8177.t182 IREF.t160 AVDD.t1472 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X846 a_n13990_8177.t181 IREF.t161 AVDD.t1473 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X847 a_5396_n6451.t4 a_n11737_n15980.t46 a_n13990_n6451.t39 AVSS.t88 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X848 AVSS.t139 AVSS.t137 AVSS.t139 AVSS.t138 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X849 a_5396_n6451.t1 a_n11737_n15980.t47 a_n13990_n6451.t38 AVSS.t85 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X850 a_n6139_n20267# a_n11737_n15980.t0 a_n11737_n15980.t1 AVSS.t178 nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X851 a_n13990_8177.t284 VP.t44 a_n13990_n6451.t97 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X852 AVDD.t649 AVDD.t648 AVDD.t649 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X853 a_n13990_8177.t180 IREF.t162 AVDD.t1474 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X854 AVDD.t647 AVDD.t646 AVDD.t647 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X855 AVDD.t645 AVDD.t644 AVDD.t645 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X856 AVDD.t643 AVDD.t642 AVDD.t643 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X857 a_5396_8177.t129 a_n11317_n20927.t1 a_5396_n6451.t31 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X858 AVDD.t641 AVDD.t640 AVDD.t641 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X859 a_n13990_8177.t179 IREF.t163 AVDD.t1475 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X860 AVDD.t639 AVDD.t637 AVDD.t639 AVDD.t638 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X861 AVDD.t636 AVDD.t635 AVDD.t636 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X862 AVDD.t634 AVDD.t633 AVDD.t634 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X863 a_n13990_n5465.t72 VN.t40 a_n13990_8177.t23 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X864 a_n13990_8177.t178 IREF.t164 AVDD.t1476 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X865 VOUT.t40 a_n11317_n20927.t1 a_5396_9163.t88 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X866 IREF.t19 IREF.t18 AVDD.t1695 AVDD.t39 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X867 AVSS.t136 AVSS.t135 AVSS.t136 AVSS.t55 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X868 a_5396_8177.t128 a_n11317_n20927.t1 a_5396_n6451.t30 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X869 VOUT.t39 a_n11317_n20927.t1 a_5396_9163.t175 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X870 AVDD.t632 AVDD.t631 AVDD.t632 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X871 AVSS.t134 AVSS.t132 AVSS.t134 AVSS.t133 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X872 AVDD.t630 AVDD.t629 AVDD.t630 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X873 a_n13990_8177.t285 VP.t45 a_n13990_n6451.t96 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X874 AVDD.t628 AVDD.t627 AVDD.t628 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X875 AVDD.t1323 a_5396_n6451.t159 a_5396_9163.t42 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X876 a_n13990_8177.t177 IREF.t165 AVDD.t1441 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X877 AVSS.t131 AVSS.t130 AVSS.t131 AVSS.t114 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X878 a_n13990_n5465.t71 VN.t41 a_n13990_8177.t24 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X879 AVDD.t626 AVDD.t625 AVDD.t626 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X880 a_5396_9163.t41 a_5396_n6451.t160 AVDD.t1324 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X881 a_5396_8177.t40 a_5396_n6451.t161 AVDD.t1325 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X882 a_n13990_8177.t25 VN.t42 a_n13990_n5465.t70 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X883 AVDD.t624 AVDD.t623 AVDD.t624 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X884 AVDD.t622 AVDD.t621 AVDD.t622 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X885 a_n13990_8177.t286 VP.t46 a_n13990_n6451.t95 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X886 AVDD.t620 AVDD.t619 AVDD.t620 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X887 VOUT.t38 a_n11317_n20927.t1 a_5396_9163.t174 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X888 AVDD.t1326 a_5396_n6451.t162 a_5396_8177.t39 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X889 AVDD.t618 AVDD.t617 AVDD.t618 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X890 a_n13990_8177.t287 VP.t47 a_n13990_n6451.t94 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X891 a_n13990_n6451.t93 VP.t48 a_n13990_8177.t73 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X892 AVDD.t1327 a_5396_n6451.t163 a_5396_9163.t40 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X893 a_n13990_8177.t176 IREF.t166 AVDD.t1442 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X894 VOUT.t37 a_n11317_n20927.t1 a_5396_9163.t109 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X895 AVDD.t1443 IREF.t167 a_n13990_8177.t175 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X896 AVDD.t616 AVDD.t615 AVDD.t616 AVDD.t131 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X897 AVDD.t614 AVDD.t613 AVDD.t614 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X898 a_5396_8177.t127 a_n11317_n20927.t1 a_5396_n6451.t33 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X899 AVDD.t612 AVDD.t611 AVDD.t612 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X900 a_n13990_8177.t26 VN.t43 a_n13990_n5465.t69 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X901 AVDD.t610 AVDD.t609 AVDD.t610 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X902 AVDD.t608 AVDD.t607 AVDD.t608 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X903 a_n13990_8177.t17 VN.t44 a_n13990_n5465.t68 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X904 AVDD.t606 AVDD.t605 AVDD.t606 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X905 AVDD.t604 AVDD.t603 AVDD.t604 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X906 AVDD.t602 AVDD.t601 AVDD.t602 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X907 AVDD.t600 AVDD.t599 AVDD.t600 AVDD.t153 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X908 a_n13990_n5465.t21 a_n11737_n14973.t63 AVSS.t332 AVSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X909 AVDD.t598 AVDD.t597 AVDD.t598 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X910 a_n13990_n5465.t10 a_n11737_n14973.t64 AVSS.t313 AVSS.t16 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X911 AVSS.t314 a_n11737_n14973.t65 a_n13990_n6451.t19 AVSS.t19 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X912 AVDD.t1444 IREF.t168 a_n11737_n14973.t16 AVDD.t638 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X913 a_n13990_n6451.t92 VP.t49 a_n13990_8177.t74 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X914 a_n13990_8177.t75 VP.t50 a_n13990_n6451.t91 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X915 AVDD.t596 AVDD.t595 AVDD.t596 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X916 a_5396_9163.t39 a_5396_n6451.t164 AVDD.t1328 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X917 AVSS.t315 a_n11737_n14973.t66 a_n13990_n5465.t11 AVSS.t201 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X918 AVDD.t594 AVDD.t593 AVDD.t594 AVDD.t153 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X919 AVDD.t592 AVDD.t591 AVDD.t592 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X920 a_n13990_8177.t174 IREF.t169 AVDD.t1445 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X921 AVDD.t1446 IREF.t170 a_n13990_8177.t173 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X922 a_n5579_n20820# a_n11737_n15980.t48 a_n6139_n20820# AVSS.t98 nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X923 AVDD.t590 AVDD.t589 AVDD.t590 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X924 a_n13990_8177.t172 IREF.t171 AVDD.t1447 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X925 a_n13990_n5465.t12 a_n11737_n14973.t67 AVSS.t316 AVSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X926 a_n13990_8177.t18 VN.t45 a_n13990_n5465.t67 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X927 a_n13990_n5465.t128 a_n11737_n15980.t49 VOUT.t95 AVSS.t67 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X928 a_5396_9163.t108 a_n11317_n20927.t1 VOUT.t36 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X929 a_n13990_n5465.t66 VN.t46 a_n13990_8177.t19 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X930 AVDD.t588 AVDD.t587 AVDD.t588 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X931 a_5396_9163.t38 a_5396_n6451.t165 AVDD.t1329 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X932 a_n13990_n5465.t127 a_n11737_n15980.t50 VOUT.t94 AVSS.t64 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X933 a_n13990_n6451.t5 a_n11737_n14973.t68 AVSS.t291 AVSS.t175 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X934 AVDD.t586 AVDD.t585 AVDD.t586 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X935 a_n13990_n5465.t65 VN.t47 a_n13990_8177.t20 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X936 a_n13990_n6451.t6 a_n11737_n14973.t69 AVSS.t292 AVSS.t172 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X937 a_5396_8177.t126 a_n11317_n20927.t1 a_5396_n6451.t32 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X938 AVSS.t129 AVSS.t128 AVSS.t129 AVSS.t74 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X939 a_5396_n6451.t31 a_n11317_n20927.t1 a_5396_8177.t125 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X940 a_n11317_n20927.t1 a_n11317_n20927.t1 a_n965_n15598# AVDD.t2 pfet_03v3 ad=0.78p pd=3.7u as=0.78p ps=3.7u w=1.2u l=2u
X941 a_n13990_8177.t21 VN.t48 a_n13990_n5465.t64 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X942 a_5396_9163.t37 a_5396_n6451.t166 AVDD.t1330 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X943 AVDD.t1448 IREF.t172 a_n13990_8177.t171 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X944 AVDD.t584 AVDD.t583 AVDD.t584 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X945 a_5396_8177.t38 a_5396_n6451.t167 AVDD.t1331 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X946 AVDD.t582 AVDD.t581 AVDD.t582 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X947 AVDD.t580 AVDD.t579 AVDD.t580 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X948 a_5396_9163.t123 a_n11317_n20927.t1 VOUT.t35 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X949 a_n13990_n5465.t63 VN.t49 a_n13990_8177.t12 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X950 AVDD.t578 AVDD.t577 AVDD.t578 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X951 AVDD.t576 AVDD.t575 AVDD.t576 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X952 a_n13990_8177.t76 VP.t51 a_n13990_n6451.t90 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X953 a_5396_n6451.t30 a_n11317_n20927.t1 a_5396_8177.t124 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X954 AVDD.t574 AVDD.t573 AVDD.t574 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X955 AVDD.t1449 IREF.t173 a_n13990_8177.t170 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X956 AVDD.t572 AVDD.t571 AVDD.t572 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X957 AVDD.t1332 a_5396_n6451.t168 a_5396_8177.t37 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X958 AVDD.t570 AVDD.t569 AVDD.t570 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X959 AVDD.t1333 a_5396_n6451.t169 a_5396_9163.t36 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X960 AVDD.t568 AVDD.t567 AVDD.t568 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X961 VOUT.t34 a_n11317_n20927.t1 a_5396_9163.t122 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X962 AVDD.t566 AVDD.t565 AVDD.t566 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X963 a_n13990_8177.t169 IREF.t174 AVDD.t1450 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X964 AVDD.t564 AVDD.t563 AVDD.t564 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X965 a_5396_8177.t123 a_n11317_n20927.t1 a_5396_n6451.t29 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X966 a_n13990_n5465.t62 VN.t50 a_n13990_8177.t13 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X967 a_n13990_n5465.t61 VN.t51 a_n13990_8177.t14 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X968 AVDD.t1451 IREF.t175 a_n13990_8177.t168 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X969 a_n13990_8177.t167 IREF.t176 AVDD.t1452 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X970 AVDD.t562 AVDD.t561 AVDD.t562 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X971 a_n13990_8177.t166 IREF.t177 AVDD.t1453 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X972 AVDD.t1454 IREF.t178 a_n13990_8177.t165 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X973 AVDD.t1334 a_5396_n6451.t170 a_5396_9163.t35 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X974 AVDD.t560 AVDD.t559 AVDD.t560 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X975 VOUT.t33 a_n11317_n20927.t1 a_5396_9163.t105 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X976 AVDD.t558 AVDD.t557 AVDD.t558 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X977 a_5396_n6451.t13 a_n11317_n20927.t1 a_5396_8177.t122 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X978 AVDD.t556 AVDD.t554 AVDD.t556 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X979 AVDD.t1335 a_5396_n6451.t171 a_5396_8177.t36 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X980 AVDD.t553 AVDD.t552 AVDD.t553 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X981 AVDD.t551 AVDD.t550 AVDD.t551 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X982 AVDD.t549 AVDD.t548 AVDD.t549 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X983 AVDD.t1336 a_5396_n6451.t172 a_5396_8177.t35 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X984 AVDD.t547 AVDD.t546 AVDD.t547 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X985 AVDD.t545 AVDD.t544 AVDD.t545 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X986 a_n11737_n14973.t15 IREF.t179 AVDD.t1455 AVDD.t39 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X987 AVDD.t543 AVDD.t542 AVDD.t543 AVDD.t2 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X988 AVSS.t127 AVSS.t126 AVSS.t127 AVSS.t49 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X989 AVDD.t541 AVDD.t540 AVDD.t541 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X990 AVDD.t539 AVDD.t538 AVDD.t539 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X991 AVDD.t1694 IREF.t16 IREF.t17 AVDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X992 AVDD.t537 AVDD.t536 AVDD.t537 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X993 a_n13990_8177.t164 IREF.t180 AVDD.t1456 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X994 AVDD.t535 AVDD.t534 AVDD.t535 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X995 AVDD.t533 AVDD.t532 AVDD.t533 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X996 AVDD.t531 AVDD.t530 AVDD.t531 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X997 a_5396_n6451.t18 a_n11317_n20927.t1 a_5396_8177.t121 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X998 AVSS.t125 AVSS.t124 AVSS.t125 AVSS.t43 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X999 AVSS.t293 a_n11737_n14973.t70 a_n13990_n6451.t7 AVSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1000 AVDD.t529 AVDD.t528 AVDD.t529 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1001 a_n13990_n6451.t89 VP.t52 a_n13990_8177.t77 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1002 AVDD.t527 AVDD.t526 AVDD.t527 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1003 AVDD.t525 AVDD.t524 AVDD.t525 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1004 AVDD.t523 AVDD.t522 AVDD.t523 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1005 AVDD.t521 AVDD.t520 AVDD.t521 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1006 AVDD.t519 AVDD.t518 AVDD.t519 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1007 a_n11737_n15980.t11 IREF.t181 AVDD.t1457 AVDD.t39 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1008 AVDD.t1693 IREF.t14 IREF.t15 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1009 a_n13990_8177.t87 VP.t53 a_n13990_n6451.t88 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1010 a_n13990_n6451.t8 a_n11737_n14973.t71 AVSS.t294 AVSS.t158 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1011 a_5396_8177.t34 a_5396_n6451.t173 AVDD.t1337 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1012 a_n13990_n6451.t21 a_n11737_n14973.t72 AVSS.t325 AVSS.t155 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1013 AVDD.t1458 IREF.t182 a_n13990_8177.t163 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1014 a_n13990_8177.t15 VN.t52 a_n13990_n5465.t60 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1015 a_5396_n6451.t61 a_n11317_n20927.t1 a_5396_8177.t120 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1016 AVDD.t1338 a_5396_n6451.t174 a_5396_8177.t33 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1017 AVDD.t517 AVDD.t516 AVDD.t517 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1018 a_n13990_8177.t16 VN.t53 a_n13990_n5465.t59 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1019 a_n13990_8177.t162 IREF.t183 AVDD.t1477 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1020 a_n13990_8177.t88 VP.t54 a_n13990_n6451.t87 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1021 AVDD.t515 AVDD.t514 AVDD.t515 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1022 a_n13990_n6451.t37 a_n11737_n15980.t51 a_5396_n6451.t3 AVSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1023 AVDD.t513 AVDD.t512 AVDD.t513 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1024 AVDD.t511 AVDD.t510 AVDD.t511 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1025 a_5396_9163.t34 a_5396_n6451.t175 AVDD.t1605 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1026 AVDD.t509 AVDD.t508 AVDD.t509 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1027 a_n13990_8177.t89 VP.t55 a_n13990_n6451.t86 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1028 AVDD.t507 AVDD.t506 AVDD.t507 AVDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1029 AVDD.t505 AVDD.t504 AVDD.t505 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1030 a_n13990_8177.t7 VN.t54 a_n13990_n5465.t58 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1031 AVDD.t503 AVDD.t502 AVDD.t503 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1032 AVDD.t501 AVDD.t500 AVDD.t501 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1033 a_5396_9163.t104 a_n11317_n20927.t1 VOUT.t32 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1034 AVDD.t1606 a_5396_n6451.t176 a_5396_8177.t32 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1035 AVDD.t499 AVDD.t498 AVDD.t499 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1036 a_5396_9163.t33 a_5396_n6451.t177 AVDD.t1607 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1037 AVDD.t497 AVDD.t496 AVDD.t497 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1038 AVDD.t495 AVDD.t494 AVDD.t495 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1039 AVDD.t1478 IREF.t184 a_n13990_8177.t161 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1040 AVDD.t1479 IREF.t185 a_n13990_8177.t160 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1041 AVDD.t1608 a_5396_n6451.t178 a_5396_8177.t31 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1042 a_n13990_8177.t159 IREF.t186 AVDD.t1480 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1043 AVDD.t1481 IREF.t187 a_n11737_n15980.t10 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1044 AVDD.t493 AVDD.t492 AVDD.t493 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1045 a_n13990_n5465.t57 VN.t55 a_n13990_8177.t8 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1046 AVSS.t123 AVSS.t122 AVSS.t123 AVSS.t55 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1047 AVDD.t491 AVDD.t490 AVDD.t491 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1048 a_n13990_8177.t90 VP.t56 a_n13990_n6451.t85 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1049 AVDD.t1482 IREF.t188 a_n13990_8177.t158 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1050 a_n13990_n5465.t18 a_n11737_n14973.t73 AVSS.t326 AVSS.t175 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1051 a_n13990_n5465.t19 a_n11737_n14973.t74 AVSS.t327 AVSS.t172 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1052 a_5396_9163.t159 a_n11317_n20927.t1 VOUT.t31 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1053 AVDD.t489 AVDD.t488 AVDD.t489 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1054 a_5396_8177.t119 a_n11317_n20927.t1 a_5396_n6451.t60 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1055 AVDD.t1609 a_5396_n6451.t179 a_5396_9163.t32 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1056 AVSS.t328 a_n11737_n14973.t75 a_n13990_n5465.t20 AVSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1057 a_n13990_n5465.t56 VN.t56 a_n13990_8177.t9 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1058 AVDD.t487 AVDD.t486 AVDD.t487 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1059 AVSS.t121 AVSS.t120 AVSS.t121 AVSS.t82 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1060 AVDD.t485 AVDD.t484 AVDD.t485 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1061 a_5396_8177.t30 a_5396_n6451.t180 AVDD.t1610 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1062 AVDD.t1611 a_5396_n6451.t181 a_5396_9163.t31 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1063 AVDD.t483 AVDD.t482 AVDD.t483 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1064 a_n13990_8177.t157 IREF.t189 AVDD.t1483 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1065 a_n13990_8177.t156 IREF.t190 AVDD.t1484 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1066 AVDD.t1485 IREF.t191 a_n13990_8177.t155 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1067 a_5396_9163.t158 a_n11317_n20927.t1 VOUT.t30 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1068 AVDD.t481 AVDD.t479 AVDD.t481 AVDD.t480 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1069 AVDD.t478 AVDD.t477 AVDD.t478 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1070 AVDD.t476 AVDD.t475 AVDD.t476 AVDD.t39 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1071 a_n11737_n14973.t14 IREF.t192 AVDD.t1486 AVDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1072 AVDD.t474 AVDD.t473 AVDD.t474 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1073 AVDD.t472 AVDD.t471 AVDD.t472 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1074 AVSS.t119 AVSS.t118 AVSS.t119 AVSS.t79 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1075 a_n13990_n6451.t84 VP.t57 a_n13990_8177.t91 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1076 AVDD.t470 AVDD.t469 AVDD.t470 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1077 AVDD.t468 AVDD.t467 AVDD.t468 AVDD.t193 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1078 a_5396_9163.t155 a_n11317_n20927.t1 VOUT.t29 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1079 a_n13990_8177.t154 IREF.t193 AVDD.t1487 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1080 AVDD.t466 AVDD.t465 AVDD.t466 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1081 AVDD.t464 AVDD.t463 AVDD.t464 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1082 AVDD.t462 AVDD.t461 AVDD.t462 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1083 AVSS.t344 a_n11737_n14973.t76 a_n13990_n6451.t29 AVSS.t235 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1084 AVDD.t460 AVDD.t459 AVDD.t460 AVDD.t193 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1085 AVDD.t458 AVDD.t457 AVDD.t458 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1086 AVDD.t456 AVDD.t455 AVDD.t456 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1087 a_5396_8177.t118 a_n11317_n20927.t1 a_5396_n6451.t59 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1088 a_5396_8177.t29 a_5396_n6451.t182 AVDD.t1612 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1089 AVDD.t1488 IREF.t194 a_n13990_8177.t153 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1090 AVDD.t1489 IREF.t195 a_n13990_8177.t152 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1091 AVDD.t454 AVDD.t453 AVDD.t454 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1092 AVDD.t452 AVDD.t451 AVDD.t452 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1093 a_5396_9163.t30 a_5396_n6451.t183 AVDD.t1613 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1094 AVSS.t117 AVSS.t116 AVSS.t117 AVSS.t25 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1095 AVSS.t345 a_n11737_n14973.t77 a_n11317_n20927.t1 AVSS.t138 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X1096 AVDD.t450 AVDD.t449 AVDD.t450 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1097 AVDD.t448 AVDD.t447 AVDD.t448 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1098 AVSS.t346 a_n11737_n14973.t78 a_n13990_n5465.t116 AVSS.t144 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1099 AVSS.t347 a_n11737_n14973.t79 a_n13990_n5465.t117 AVSS.t141 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1100 AVDD.t446 AVDD.t445 AVDD.t446 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1101 a_n13990_n6451.t83 VP.t58 a_n13990_8177.t63 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1102 a_n13990_n6451.t82 VP.t59 a_n13990_8177.t64 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1103 AVDD.t1490 IREF.t196 a_n13990_8177.t151 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1104 AVDD.t444 AVDD.t443 AVDD.t444 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1105 a_n13990_n6451.t81 VP.t60 a_n13990_8177.t65 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1106 AVDD.t1614 a_5396_n6451.t184 a_5396_8177.t28 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1107 AVDD.t442 AVDD.t441 AVDD.t442 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1108 AVDD.t440 AVDD.t439 AVDD.t440 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1109 a_5396_n6451.t39 a_n11317_n20927.t1 a_5396_8177.t117 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1110 AVDD.t438 AVDD.t437 AVDD.t438 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1111 AVDD.t1491 IREF.t197 a_n13990_8177.t150 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1112 AVDD.t436 AVDD.t435 AVDD.t436 AVDD.t2 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1113 VOUT.t28 a_n11317_n20927.t1 a_5396_9163.t154 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1114 a_5396_n6451.t58 a_n11317_n20927.t1 a_5396_8177.t116 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1115 VOUT.t93 a_n11737_n15980.t52 a_n13990_n5465.t138 AVSS.t88 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1116 VOUT.t92 a_n11737_n15980.t53 a_n13990_n5465.t137 AVSS.t85 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1117 a_n13990_n6451.t80 VP.t61 a_n13990_8177.t66 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1118 a_5396_n6451.t26 a_n11317_n20927.t1 a_5396_8177.t115 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1119 AVDD.t434 AVDD.t433 AVDD.t434 AVDD.t178 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1120 AVDD.t432 AVDD.t431 AVDD.t432 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1121 AVSS.t115 AVSS.t113 AVSS.t115 AVSS.t114 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1122 AVDD.t430 AVDD.t429 AVDD.t430 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1123 AVDD.t1492 IREF.t198 a_n13990_8177.t149 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1124 AVSS.t352 a_n11737_n14973.t0 a_n11737_n14973.t1 AVSS.t133 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X1125 AVDD.t1615 a_5396_n6451.t185 a_5396_8177.t27 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1126 AVDD.t428 AVDD.t427 AVDD.t428 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1127 a_5396_8177.t114 a_n11317_n20927.t1 a_5396_n6451.t22 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1128 AVSS.t112 AVSS.t111 AVSS.t112 AVSS.t49 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1129 AVDD.t426 AVDD.t425 AVDD.t426 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1130 AVDD.t1493 IREF.t199 a_n13990_8177.t148 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1131 a_n13990_8177.t147 IREF.t200 AVDD.t1494 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1132 AVDD.t424 AVDD.t423 AVDD.t424 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1133 AVDD.t422 AVDD.t421 AVDD.t422 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1134 VOUT.t27 a_n11317_n20927.t5 a_5396_9163.t153 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1135 VOUT.t26 a_n11317_n20927.t1 a_5396_9163.t152 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1136 a_n11737_n15980.t9 IREF.t201 AVDD.t1380 AVDD.t480 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1137 a_n13990_n5465.t7 a_n11737_n14973.t80 AVSS.t309 AVSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1138 AVDD.t420 AVDD.t419 AVDD.t420 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1139 AVDD.t1381 IREF.t202 a_n11737_n14973.t13 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1140 AVDD.t1616 a_5396_n6451.t186 a_5396_9163.t29 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1141 AVDD.t418 AVDD.t417 AVDD.t418 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1142 a_5396_9163.t145 a_n11317_n20927.t1 VOUT.t25 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1143 AVDD.t416 AVDD.t415 AVDD.t416 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1144 a_n13990_n5465.t8 a_n11737_n14973.t81 AVSS.t310 AVSS.t158 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1145 a_n13990_8177.t67 VP.t62 a_n13990_n6451.t79 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1146 a_n13990_n5465.t9 a_n11737_n14973.t82 AVSS.t311 AVSS.t155 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1147 a_n13990_n6451.t18 a_n11737_n14973.t83 AVSS.t312 AVSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1148 AVDD.t1617 a_5396_n6451.t187 a_5396_9163.t28 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1149 AVSS.t287 a_n11737_n14973.t84 a_n13990_n5465.t1 AVSS.t19 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1150 a_n13990_n6451.t3 a_n11737_n14973.t85 AVSS.t288 AVSS.t16 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1151 AVDD.t414 AVDD.t413 AVDD.t414 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1152 AVDD.t412 AVDD.t411 AVDD.t412 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1153 VOUT.t91 a_n11737_n15980.t54 a_n13990_n5465.t134 AVSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1154 VOUT.t24 a_n11317_n20927.t1 a_5396_9163.t144 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1155 AVDD.t1382 IREF.t203 a_n11737_n14973.t12 AVDD.t810 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1156 VOUT.t90 a_n11737_n15980.t55 a_n13990_n5465.t133 AVSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1157 AVDD.t410 AVDD.t409 AVDD.t410 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1158 a_n13990_8177.t10 VN.t57 a_n13990_n5465.t55 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1159 AVDD.t1383 IREF.t204 a_n13990_8177.t146 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1160 AVDD.t1384 IREF.t205 a_n11737_n15980.t8 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1161 AVDD.t408 AVDD.t407 AVDD.t408 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1162 AVDD.t1618 a_5396_n6451.t188 a_5396_8177.t26 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1163 a_5396_9163.t27 a_5396_n6451.t189 AVDD.t1619 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1164 a_5396_8177.t113 a_n11317_n20927.t1 a_5396_n6451.t53 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1165 AVDD.t1620 a_5396_n6451.t190 a_5396_9163.t26 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1166 AVDD.t406 AVDD.t405 AVDD.t406 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1167 AVDD.t404 AVDD.t403 AVDD.t404 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1168 AVDD.t1385 IREF.t206 a_n13990_8177.t145 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1169 AVSS.t110 AVSS.t109 AVSS.t110 AVSS.t98 nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X1170 AVDD.t402 AVDD.t401 AVDD.t402 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1171 AVDD.t400 AVDD.t398 AVDD.t400 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1172 a_n13990_8177.t11 VN.t58 a_n13990_n5465.t54 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1173 a_5396_8177.t25 a_5396_n6451.t191 AVDD.t1621 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1174 AVDD.t397 AVDD.t396 AVDD.t397 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1175 a_n13990_8177.t144 IREF.t207 AVDD.t1386 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1176 AVDD.t395 AVDD.t393 AVDD.t395 AVDD.t394 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X1177 AVDD.t392 AVDD.t391 AVDD.t392 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1178 AVSS.t289 a_n11737_n14973.t86 a_n13990_n5465.t2 AVSS.t222 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1179 AVDD.t390 AVDD.t389 AVDD.t390 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1180 a_5396_8177.t24 a_5396_n6451.t192 AVDD.t1622 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1181 AVDD.t388 AVDD.t387 AVDD.t388 AVDD.t13 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1182 AVDD.t386 AVDD.t385 AVDD.t386 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1183 AVDD.t1387 IREF.t208 a_n13990_8177.t143 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1184 AVDD.t1388 IREF.t209 a_n13990_8177.t142 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1185 a_n13990_n6451.t36 a_n11737_n15980.t56 a_5396_n6451.t2 AVSS.t67 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1186 AVDD.t384 AVDD.t383 AVDD.t384 AVDD.t156 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1187 a_n13990_n6451.t35 a_n11737_n15980.t57 a_5396_n6451.t63 AVSS.t64 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1188 AVDD.t382 AVDD.t380 AVDD.t382 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1189 a_n13990_n6451.t78 VP.t63 a_n13990_8177.t322 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1190 AVDD.t379 AVDD.t377 AVDD.t379 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1191 AVDD.t376 AVDD.t375 AVDD.t376 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1192 a_n13990_8177.t141 IREF.t210 AVDD.t1389 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1193 a_n13990_8177.t323 VP.t64 a_n13990_n6451.t77 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1194 a_5396_8177.t23 a_5396_n6451.t193 AVDD.t1623 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1195 AVDD.t1624 a_5396_n6451.t194 a_5396_9163.t25 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1196 AVDD.t1625 a_5396_n6451.t195 a_5396_8177.t22 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1197 a_n11737_n15980.t7 IREF.t211 AVDD.t1390 AVDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1198 AVDD.t1391 IREF.t212 a_n13990_8177.t140 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1199 a_5396_8177.t112 a_n11317_n20927.t1 a_5396_n6451.t57 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1200 AVDD.t374 AVDD.t372 AVDD.t374 AVDD.t373 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1201 AVSS.t108 AVSS.t107 AVSS.t108 AVSS.t74 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1202 a_5396_8177.t111 a_n11317_n20927.t1 a_5396_n6451.t56 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1203 a_5396_8177.t110 a_n11317_n20927.t1 a_5396_n6451.t55 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1204 a_n13990_8177.t324 VP.t65 a_n13990_n6451.t76 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1205 VOUT.t23 a_n11317_n20927.t1 a_5396_9163.t97 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1206 a_5396_9163.t96 a_n11317_n20927.t1 VOUT.t22 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1207 a_n13990_8177.t139 IREF.t213 AVDD.t1392 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1208 AVDD.t371 AVDD.t370 AVDD.t371 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1209 AVDD.t369 AVDD.t368 AVDD.t369 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1210 AVDD.t367 AVDD.t365 AVDD.t367 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1211 AVSS.t106 AVSS.t105 AVSS.t106 AVSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1212 AVDD.t364 AVDD.t363 AVDD.t364 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1213 AVDD.t362 AVDD.t361 AVDD.t362 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1214 a_n13990_n6451.t4 a_n11737_n14973.t87 AVSS.t290 AVSS.t144 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1215 AVSS.t104 AVSS.t102 AVSS.t104 AVSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1216 a_n13990_n6451.t49 a_n11737_n14973.t88 AVSS.t354 AVSS.t141 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1217 a_n13990_8177.t138 IREF.t214 AVDD.t1393 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1218 AVSS.t101 AVSS.t100 AVSS.t101 AVSS.t1 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1219 AVDD.t360 AVDD.t359 AVDD.t360 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1220 a_n13990_8177.t137 IREF.t215 AVDD.t1394 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1221 AVDD.t358 AVDD.t357 AVDD.t358 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1222 AVSS.t99 AVSS.t97 AVSS.t99 AVSS.t98 nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X1223 a_5396_9163.t151 a_n11317_n20927.t1 VOUT.t21 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1224 a_n13990_8177.t325 VP.t66 a_n13990_n6451.t75 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1225 a_n13990_n5465.t53 VN.t59 a_n13990_8177.t82 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1226 AVDD.t1395 IREF.t216 a_n13990_8177.t136 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1227 AVSS.t96 AVSS.t94 AVSS.t96 AVSS.t95 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X1228 VOUT.t20 a_n11317_n20927.t1 a_5396_9163.t150 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1229 a_5396_9163.t24 a_5396_n6451.t196 AVDD.t1626 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1230 AVDD.t356 AVDD.t355 AVDD.t356 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1231 AVDD.t354 AVDD.t353 AVDD.t354 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1232 a_5396_8177.t109 a_n11317_n20927.t1 a_5396_n6451.t28 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1233 AVDD.t1396 IREF.t217 a_n13990_8177.t135 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1234 a_5396_8177.t108 a_n11317_n20927.t1 a_5396_n6451.t14 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1235 AVDD.t1627 a_5396_n6451.t197 a_5396_9163.t23 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1236 VOUT.t89 a_n11737_n15980.t58 a_n13990_n5465.t124 AVSS.t37 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1237 AVSS.t93 AVSS.t92 AVSS.t93 AVSS.t43 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1238 a_5396_9163.t125 a_n11317_n20927.t1 VOUT.t19 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1239 AVDD.t352 AVDD.t351 AVDD.t352 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1240 a_n13990_n5465.t52 VN.t60 a_n13990_8177.t83 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1241 AVDD.t1628 a_5396_n6451.t198 a_5396_9163.t22 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1242 AVDD.t1629 a_5396_n6451.t199 a_5396_8177.t21 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1243 AVDD.t350 AVDD.t349 AVDD.t350 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1244 a_n13990_n6451.t74 VP.t67 a_n13990_8177.t326 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1245 AVDD.t348 AVDD.t346 AVDD.t348 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1246 a_5396_n6451.t51 a_n11317_n20927.t1 a_5396_8177.t107 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1247 AVDD.t345 AVDD.t344 AVDD.t345 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1248 AVDD.t1397 IREF.t218 a_n13990_8177.t134 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1249 AVDD.t343 AVDD.t342 AVDD.t343 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1250 AVDD.t341 AVDD.t340 AVDD.t341 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1251 AVDD.t339 AVDD.t337 AVDD.t339 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1252 AVDD.t336 AVDD.t334 AVDD.t336 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1253 a_5396_9163.t21 a_5396_n6451.t200 AVDD.t1630 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1254 a_5396_9163.t20 a_5396_n6451.t201 AVDD.t1631 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1255 AVDD.t333 AVDD.t332 AVDD.t333 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1256 a_5396_9163.t124 a_n11317_n20927.t1 VOUT.t18 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1257 a_n13990_8177.t133 IREF.t219 AVDD.t1398 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1258 AVSS.t91 AVSS.t90 AVSS.t91 AVSS.t34 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1259 a_5396_n6451.t54 a_n11317_n20927.t1 a_5396_8177.t106 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1260 a_n13990_8177.t132 IREF.t220 AVDD.t1399 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1261 a_n13990_8177.t131 IREF.t221 AVDD.t1400 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1262 a_n13990_8177.t84 VN.t61 a_n13990_n5465.t51 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1263 IREF.t13 IREF.t12 AVDD.t1692 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1264 AVSS.t355 a_n11737_n14973.t89 a_n13990_n6451.t50 AVSS.t201 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1265 AVDD.t331 AVDD.t330 AVDD.t331 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1266 AVDD.t329 AVDD.t327 AVDD.t329 AVDD.t328 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1267 a_n13990_8177.t130 IREF.t222 AVDD.t1401 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1268 AVDD.t326 AVDD.t325 AVDD.t326 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1269 a_n13990_n6451.t73 VP.t68 a_n13990_8177.t312 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1270 a_5396_8177.t20 a_5396_n6451.t202 AVDD.t1632 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1271 IREF.t11 IREF.t10 AVDD.t1691 AVDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1272 AVDD.t324 AVDD.t322 AVDD.t324 AVDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1273 a_5396_9163.t19 a_5396_n6451.t203 AVDD.t1633 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1274 a_n13990_n6451.t72 VP.t69 a_n13990_8177.t313 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1275 AVDD.t1634 a_5396_n6451.t204 a_5396_8177.t19 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1276 a_5396_n6451.t54 a_n11317_n20927.t1 a_5396_8177.t105 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1277 AVDD.t321 AVDD.t320 AVDD.t321 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1278 a_n13990_8177.t85 VN.t62 a_n13990_n5465.t50 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1279 AVDD.t319 AVDD.t318 AVDD.t319 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1280 AVDD.t317 AVDD.t316 AVDD.t317 AVDD.t156 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1281 a_n13990_8177.t129 IREF.t223 AVDD.t1402 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1282 AVDD.t315 AVDD.t314 AVDD.t315 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1283 AVDD.t313 AVDD.t312 AVDD.t313 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1284 AVDD.t1635 a_5396_n6451.t205 a_5396_9163.t18 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1285 a_5396_9163.t17 a_5396_n6451.t206 AVDD.t1636 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1286 AVDD.t311 AVDD.t310 AVDD.t311 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1287 a_n13990_8177.t314 VP.t70 a_n13990_n6451.t71 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1288 AVDD.t309 AVDD.t308 AVDD.t309 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1289 a_5396_8177.t104 a_n11317_n20927.t1 a_5396_n6451.t48 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1290 AVDD.t1637 a_5396_n6451.t207 a_5396_9163.t16 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1291 AVSS.t89 AVSS.t87 AVSS.t89 AVSS.t88 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1292 AVSS.t86 AVSS.t84 AVSS.t86 AVSS.t85 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1293 AVSS.t83 AVSS.t81 AVSS.t83 AVSS.t82 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1294 AVDD.t1638 a_5396_n6451.t208 a_5396_8177.t18 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1295 AVDD.t307 AVDD.t306 AVDD.t307 AVDD.t193 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1296 AVSS.t356 a_n11737_n14973.t90 a_n13990_n5465.t139 AVSS.t235 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1297 AVDD.t305 AVDD.t304 AVDD.t305 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1298 AVDD.t1403 IREF.t224 a_n13990_8177.t128 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1299 AVDD.t303 AVDD.t302 AVDD.t303 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1300 a_n13990_8177.t315 VP.t71 a_n13990_n6451.t70 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1301 a_n13990_8177.t316 VP.t72 a_n13990_n6451.t69 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1302 AVSS.t80 AVSS.t78 AVSS.t80 AVSS.t79 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1303 AVDD.t1639 a_5396_n6451.t209 a_5396_9163.t15 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1304 AVDD.t301 AVDD.t300 AVDD.t301 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1305 a_n13990_n6451.t34 a_n11737_n15980.t59 a_5396_n6451.t0 AVSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1306 a_5396_n6451.t28 a_n11317_n20927.t1 a_5396_8177.t103 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1307 AVDD.t299 AVDD.t298 AVDD.t299 AVDD.t156 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1308 a_n13990_8177.t86 VN.t63 a_n13990_n5465.t49 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1309 a_5396_8177.t17 a_5396_n6451.t210 AVDD.t1495 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1310 a_n13990_n6451.t68 VP.t73 a_n13990_8177.t48 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1311 a_5396_9163.t14 a_5396_n6451.t211 AVDD.t1496 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1312 a_n13990_8177.t127 IREF.t225 AVDD.t1404 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1313 a_n13990_8177.t342 VN.t64 a_n13990_n5465.t48 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1314 AVSS.t77 AVSS.t76 AVSS.t77 AVSS.t25 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1315 a_5396_9163.t135 a_n11317_n20927.t1 VOUT.t17 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1316 AVDD.t297 AVDD.t296 AVDD.t297 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1317 AVDD.t295 AVDD.t293 AVDD.t295 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1318 AVSS.t75 AVSS.t73 AVSS.t75 AVSS.t74 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1319 a_n13990_8177.t126 IREF.t226 AVDD.t1405 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1320 AVDD.t292 AVDD.t290 AVDD.t292 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1321 a_5396_9163.t134 a_n11317_n20927.t1 VOUT.t16 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1322 AVDD.t1406 IREF.t227 a_n13990_8177.t125 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1323 a_n13990_8177.t343 VN.t65 a_n13990_n5465.t47 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1324 a_5396_n6451.t25 a_n11317_n20927.t1 a_5396_8177.t102 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1325 AVDD.t289 AVDD.t288 AVDD.t289 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1326 a_n11737_n15980.t6 IREF.t228 AVDD.t1407 AVDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1327 a_n13990_8177.t344 VN.t66 a_n13990_n5465.t46 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1328 AVDD.t1497 a_5396_n6451.t212 a_5396_9163.t13 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1329 AVDD.t1498 a_5396_n6451.t213 a_5396_8177.t16 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1330 AVDD.t1499 a_5396_n6451.t214 a_5396_9163.t12 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1331 AVDD.t287 AVDD.t286 AVDD.t287 AVDD.t153 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1332 AVDD.t285 AVDD.t284 AVDD.t285 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1333 AVDD.t283 AVDD.t281 AVDD.t283 AVDD.t282 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1334 a_5396_9163.t133 a_n11317_n20927.t1 VOUT.t15 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1335 a_5396_8177.t101 a_n11317_n20927.t1 a_5396_n6451.t27 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1336 AVDD.t280 AVDD.t278 AVDD.t280 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1337 AVDD.t277 AVDD.t276 AVDD.t277 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1338 AVSS.t72 AVSS.t71 AVSS.t72 AVSS.t46 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1339 a_5396_9163.t132 a_n11317_n20927.t1 VOUT.t14 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1340 AVDD.t1285 IREF.t8 IREF.t9 AVDD.t810 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1341 AVDD.t275 AVDD.t274 AVDD.t275 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1342 a_n13990_8177.t345 VN.t67 a_n13990_n5465.t45 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1343 AVDD.t273 AVDD.t272 AVDD.t273 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1344 a_5396_8177.t100 a_n11317_n20927.t1 a_5396_n6451.t26 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1345 a_5396_n6451.t25 a_n11317_n20927.t1 a_5396_8177.t99 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1346 a_n13990_8177.t346 VN.t68 a_n13990_n5465.t44 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1347 AVDD.t1284 IREF.t6 IREF.t7 AVDD.t638 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1348 AVDD.t271 AVDD.t270 AVDD.t271 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1349 AVDD.t269 AVDD.t268 AVDD.t269 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1350 AVDD.t267 AVDD.t266 AVDD.t267 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1351 AVDD.t265 AVDD.t263 AVDD.t265 AVDD.t264 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X1352 AVDD.t262 AVDD.t261 AVDD.t262 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1353 a_5396_9163.t121 a_n11317_n20927.t1 VOUT.t13 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1354 a_n13990_n6451.t33 a_n11737_n15980.t60 a_5396_n6451.t1 AVSS.t37 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1355 a_n13990_n5465.t43 VN.t69 a_n13990_8177.t53 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1356 a_n13990_8177.t124 IREF.t229 AVDD.t1408 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1357 AVDD.t260 AVDD.t259 AVDD.t260 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1358 a_n13990_8177.t54 VN.t70 a_n13990_n5465.t42 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1359 AVDD.t258 AVDD.t257 AVDD.t258 AVDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1360 AVDD.t256 AVDD.t254 AVDD.t256 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1361 a_5396_9163.t120 a_n11317_n20927.t1 VOUT.t12 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1362 AVDD.t253 AVDD.t251 AVDD.t253 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1363 a_n13990_n5465.t41 VN.t71 a_n13990_8177.t55 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1364 a_n13990_8177.t123 IREF.t230 AVDD.t1409 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1365 AVSS.t70 AVSS.t69 AVSS.t70 AVSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1366 a_5396_9163.t11 a_5396_n6451.t215 AVDD.t1500 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1367 AVSS.t68 AVSS.t66 AVSS.t68 AVSS.t67 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1368 AVDD.t250 AVDD.t249 AVDD.t250 AVDD.t178 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1369 a_5396_8177.t15 a_5396_n6451.t216 AVDD.t1501 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1370 a_5396_8177.t14 a_5396_n6451.t217 AVDD.t1502 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1371 AVSS.t65 AVSS.t63 AVSS.t65 AVSS.t64 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1372 AVDD.t248 AVDD.t247 AVDD.t248 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1373 a_5396_9163.t171 a_n11317_n20927.t1 VOUT.t11 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1374 AVDD.t1410 IREF.t231 a_n13990_8177.t122 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1375 AVDD.t246 AVDD.t245 AVDD.t246 AVDD.t181 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1376 a_n13990_n6451.t51 a_n11737_n14973.t91 AVSS.t357 AVSS.t114 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1377 AVDD.t244 AVDD.t243 AVDD.t244 AVDD.t178 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1378 AVDD.t242 AVDD.t240 AVDD.t242 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1379 AVDD.t239 AVDD.t237 AVDD.t239 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1380 a_n13990_n6451.t67 VP.t74 a_n13990_8177.t49 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1381 AVDD.t236 AVDD.t235 AVDD.t236 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1382 a_5396_8177.t98 a_n11317_n20927.t1 a_5396_n6451.t24 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1383 AVDD.t234 AVDD.t232 AVDD.t234 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1384 AVSS.t62 AVSS.t61 AVSS.t62 AVSS.t1 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1385 AVSS.t60 AVSS.t59 AVSS.t60 AVSS.t34 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1386 AVDD.t1503 a_5396_n6451.t218 a_5396_9163.t10 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1387 AVDD.t231 AVDD.t230 AVDD.t231 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1388 AVDD.t229 AVDD.t228 AVDD.t229 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1389 a_n13990_n5465.t40 VN.t72 a_n13990_8177.t56 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1390 AVDD.t227 AVDD.t225 AVDD.t227 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1391 AVDD.t224 AVDD.t223 AVDD.t224 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1392 AVDD.t222 AVDD.t221 AVDD.t222 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1393 a_n13990_n5465.t39 VN.t73 a_n13990_8177.t57 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1394 a_n13990_n6451.t15 a_n11737_n14973.t92 AVSS.t305 AVSS.t175 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1395 a_n13990_n6451.t16 a_n11737_n14973.t93 AVSS.t306 AVSS.t172 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1396 AVDD.t220 AVDD.t219 AVDD.t220 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1397 a_n13990_8177.t121 IREF.t232 AVDD.t1411 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1398 AVDD.t1412 IREF.t233 a_n11737_n15980.t5 AVDD.t282 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1399 AVDD.t218 AVDD.t217 AVDD.t218 AVDD.t193 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1400 a_n13990_n5465.t38 VN.t74 a_n13990_8177.t2 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1401 a_5396_8177.t13 a_5396_n6451.t219 AVDD.t1504 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1402 AVDD.t216 AVDD.t215 AVDD.t216 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1403 a_5396_n6451.t63 a_n11737_n15980.t61 a_n13990_n6451.t32 AVSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1404 a_5396_n6451.t3 a_n11737_n15980.t62 a_n13990_n6451.t31 AVSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1405 VOUT.t10 a_n11317_n20927.t1 a_5396_9163.t170 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1406 AVSS.t307 a_n11737_n14973.t94 a_n13990_n6451.t17 AVSS.t222 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1407 a_n13990_8177.t50 VP.t75 a_n13990_n6451.t66 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1408 AVSS.t58 AVSS.t57 AVSS.t58 AVSS.t28 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1409 AVDD.t1427 IREF.t234 a_n11737_n15980.t4 AVDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1410 AVDD.t214 AVDD.t213 AVDD.t214 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1411 a_n13990_n5465.t37 VN.t75 a_n13990_8177.t3 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1412 AVDD.t212 AVDD.t211 AVDD.t212 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1413 a_n5579_n20820# a_n11737_n15980.t63 a_n6139_n20267# AVSS.t98 nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X1414 a_5396_8177.t12 a_5396_n6451.t220 AVDD.t1505 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1415 AVDD.t210 AVDD.t209 AVDD.t210 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1416 a_5396_9163.t99 a_n11317_n20927.t1 VOUT.t9 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1417 a_n13990_n5465.t36 VN.t76 a_n13990_8177.t4 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1418 a_5396_8177.t11 a_5396_n6451.t221 AVDD.t1506 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1419 a_5396_9163.t9 a_5396_n6451.t222 AVDD.t1507 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1420 AVDD.t208 AVDD.t207 AVDD.t208 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1421 AVDD.t206 AVDD.t204 AVDD.t206 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1422 AVDD.t203 AVDD.t202 AVDD.t203 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1423 a_n1533_n16909# a_n11317_n20927.t1 a_n2101_n16909# AVDD.t394 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X1424 AVDD.t201 AVDD.t199 AVDD.t201 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1425 AVDD.t1428 IREF.t235 a_n13990_8177.t120 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1426 a_n13990_8177.t119 IREF.t236 AVDD.t1429 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1427 AVDD.t1430 IREF.t237 a_n13990_8177.t118 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1428 a_5396_8177.t10 a_5396_n6451.t223 AVDD.t1508 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1429 AVDD.t198 AVDD.t197 AVDD.t198 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1430 AVDD.t196 AVDD.t195 AVDD.t196 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1431 a_5396_8177.t9 a_5396_n6451.t224 AVDD.t1509 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1432 AVDD.t194 AVDD.t192 AVDD.t194 AVDD.t193 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1433 AVDD.t191 AVDD.t190 AVDD.t191 AVDD.t131 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1434 a_n13990_8177.t51 VP.t76 a_n13990_n6451.t65 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1435 AVDD.t189 AVDD.t188 AVDD.t189 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1436 AVDD.t187 AVDD.t185 AVDD.t187 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1437 a_5396_9163.t98 a_n11317_n20927.t1 VOUT.t8 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1438 AVDD.t184 AVDD.t183 AVDD.t184 AVDD.t153 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1439 AVDD.t182 AVDD.t180 AVDD.t182 AVDD.t181 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1440 AVSS.t56 AVSS.t54 AVSS.t56 AVSS.t55 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1441 VOUT.t7 a_n11317_n20927.t1 a_5396_9163.t95 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1442 VOUT.t88 a_n11737_n15980.t64 a_n13990_n5465.t123 AVSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1443 a_n13990_8177.t117 IREF.t238 AVDD.t1431 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1444 a_n13990_8177.t116 IREF.t239 AVDD.t1432 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1445 a_n13990_n5465.t35 VN.t77 a_n13990_8177.t5 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1446 AVDD.t1510 a_5396_n6451.t225 a_5396_9163.t8 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1447 a_n13990_n6451.t64 VP.t77 a_n13990_8177.t52 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1448 AVDD.t179 AVDD.t177 AVDD.t179 AVDD.t178 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1449 AVSS.t53 AVSS.t51 AVSS.t53 AVSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1450 AVDD.t176 AVDD.t174 AVDD.t176 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1451 AVDD.t173 AVDD.t172 AVDD.t173 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1452 AVDD.t1511 a_5396_n6451.t226 a_5396_8177.t8 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1453 AVDD.t171 AVDD.t170 AVDD.t171 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1454 AVDD.t169 AVDD.t168 AVDD.t169 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1455 AVDD.t167 AVDD.t166 AVDD.t167 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1456 VOUT.t6 a_n11317_n20927.t1 a_5396_9163.t94 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1457 AVSS.t50 AVSS.t48 AVSS.t50 AVSS.t49 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1458 a_n13990_n5465.t34 VN.t78 a_n13990_8177.t6 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1459 AVDD.t165 AVDD.t164 AVDD.t165 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1460 AVDD.t163 AVDD.t162 AVDD.t163 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1461 AVDD.t161 AVDD.t160 AVDD.t161 AVDD.t156 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1462 a_5396_8177.t7 a_5396_n6451.t227 AVDD.t1512 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1463 a_n13990_n6451.t63 VP.t78 a_n13990_8177.t68 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1464 a_5396_8177.t97 a_n11317_n20927.t1 a_5396_n6451.t23 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1465 AVDD.t159 AVDD.t158 AVDD.t159 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1466 a_n13990_8177.t115 IREF.t240 AVDD.t1433 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1467 AVDD.t1434 IREF.t241 a_n11737_n15980.t3 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1468 a_n11317_n20927.t0 a_n11737_n14973.t95 AVSS.t308 AVSS.t95 nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X1469 a_5396_9163.t149 a_n11317_n20927.t1 VOUT.t5 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1470 AVDD.t157 AVDD.t155 AVDD.t157 AVDD.t156 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1471 AVDD.t154 AVDD.t152 AVDD.t154 AVDD.t153 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1472 AVDD.t151 AVDD.t150 AVDD.t151 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1473 a_n13990_n6451.t0 a_n11737_n14973.t96 AVSS.t283 AVSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1474 AVDD.t149 AVDD.t147 AVDD.t149 AVDD.t148 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1475 AVDD.t1435 IREF.t242 a_n13990_8177.t114 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1476 AVDD.t146 AVDD.t145 AVDD.t146 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1477 a_5396_n6451.t22 a_n11317_n20927.t1 a_5396_8177.t96 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1478 a_n13990_8177.t69 VP.t79 a_n13990_n6451.t62 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1479 AVDD.t144 AVDD.t143 AVDD.t144 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1480 AVDD.t1436 IREF.t243 a_n11737_n14973.t11 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1481 AVDD.t142 AVDD.t140 AVDD.t142 AVDD.t141 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1482 a_5396_8177.t6 a_5396_n6451.t228 AVDD.t1513 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1483 a_n13990_n6451.t1 a_n11737_n14973.t97 AVSS.t284 AVSS.t158 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1484 a_n13990_n6451.t2 a_n11737_n14973.t98 AVSS.t285 AVSS.t155 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1485 a_5396_9163.t148 a_n11317_n20927.t1 VOUT.t4 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1486 AVDD.t139 AVDD.t138 AVDD.t139 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1487 IREF.t5 IREF.t4 AVDD.t1283 AVDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1488 a_5396_8177.t5 a_5396_n6451.t229 AVDD.t1514 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1489 AVDD.t137 AVDD.t135 AVDD.t137 AVDD.t136 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1490 AVSS.t286 a_n11737_n14973.t99 a_n13990_n5465.t0 AVSS.t201 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1491 a_n13990_n6451.t61 VP.t80 a_n13990_8177.t70 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1492 AVDD.t134 AVDD.t133 AVDD.t134 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1493 a_5396_9163.t7 a_5396_n6451.t230 AVDD.t1515 AVDD.t156 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1494 AVDD.t132 AVDD.t130 AVDD.t132 AVDD.t131 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1495 AVSS.t47 AVSS.t45 AVSS.t47 AVSS.t46 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1496 a_5396_n6451.t21 a_n11317_n20927.t1 a_5396_8177.t95 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1497 a_n13990_n6451.t60 VP.t81 a_n13990_8177.t71 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1498 a_5396_n6451.t44 a_n11317_n20927.t1 a_5396_8177.t94 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1499 AVDD.t129 AVDD.t128 AVDD.t129 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1500 AVSS.t44 AVSS.t42 AVSS.t44 AVSS.t43 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1501 AVSS.t340 a_n11737_n14973.t100 a_n13990_n5465.t113 AVSS.t114 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1502 a_n2101_n16909# a_n11317_n20927.t1 a_n2631_n17634# AVDD.t328 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X1503 a_n13990_n5465.t33 VN.t79 a_n13990_8177.t332 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1504 a_5396_9163.t119 a_n11317_n20927.t1 VOUT.t3 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1505 a_n13990_n6451.t59 VP.t82 a_n13990_8177.t72 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1506 AVSS.t41 AVSS.t39 AVSS.t41 AVSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1507 a_n13990_8177.t113 IREF.t244 AVDD.t1437 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1508 a_n13990_8177.t333 VN.t80 a_n13990_n5465.t32 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1509 a_5396_n6451.t21 a_n11317_n20927.t1 a_5396_8177.t93 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1510 a_n13990_n6451.t58 VP.t83 a_n13990_8177.t58 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1511 AVDD.t1438 IREF.t245 a_n13990_8177.t112 AVDD.t153 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1512 AVDD.t127 AVDD.t126 AVDD.t127 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1513 a_n13990_8177.t59 VP.t84 a_n13990_n6451.t57 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1514 AVDD.t125 AVDD.t124 AVDD.t125 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1515 a_5396_9163.t6 a_5396_n6451.t231 AVDD.t1516 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1516 AVDD.t123 AVDD.t121 AVDD.t123 AVDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1517 AVDD.t120 AVDD.t118 AVDD.t120 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1518 a_5396_9163.t5 a_5396_n6451.t232 AVDD.t1517 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1519 a_n13990_n5465.t31 VN.t81 a_n13990_8177.t334 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1520 a_n13990_8177.t335 VN.t82 a_n13990_n5465.t30 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1521 AVDD.t1439 IREF.t246 a_n13990_8177.t111 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1522 AVDD.t117 AVDD.t116 AVDD.t117 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1523 AVDD.t115 AVDD.t113 AVDD.t115 AVDD.t114 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1524 AVDD.t1282 IREF.t2 IREF.t3 AVDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1525 AVSS.t38 AVSS.t36 AVSS.t38 AVSS.t37 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1526 AVDD.t112 AVDD.t110 AVDD.t112 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1527 AVDD.t109 AVDD.t108 AVDD.t109 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1528 AVDD.t107 AVDD.t106 AVDD.t107 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1529 AVDD.t105 AVDD.t104 AVDD.t105 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1530 AVDD.t103 AVDD.t102 AVDD.t103 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1531 a_n13990_8177.t110 IREF.t247 AVDD.t1440 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1532 AVDD.t1413 IREF.t248 a_n13990_8177.t109 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1533 a_n13990_n6451.t56 VP.t85 a_n13990_8177.t60 AVDD.t294 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1534 AVDD.t101 AVDD.t100 AVDD.t101 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1535 AVDD.t99 AVDD.t97 AVDD.t99 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1536 AVDD.t96 AVDD.t95 AVDD.t96 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1537 AVDD.t94 AVDD.t92 AVDD.t94 AVDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1538 AVDD.t91 AVDD.t90 AVDD.t91 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1539 AVDD.t89 AVDD.t87 AVDD.t89 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1540 AVDD.t86 AVDD.t84 AVDD.t86 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1541 a_n11737_n15980.t2 IREF.t249 AVDD.t1414 AVDD.t638 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1542 a_n13990_n6451.t55 VP.t86 a_n13990_8177.t61 AVDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1543 AVDD.t83 AVDD.t81 AVDD.t83 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1544 a_n11737_n14973.t10 IREF.t250 AVDD.t1415 AVDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1545 AVDD.t80 AVDD.t78 AVDD.t80 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1546 AVDD.t77 AVDD.t76 AVDD.t77 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1547 AVDD.t75 AVDD.t74 AVDD.t75 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1548 AVDD.t1518 a_5396_n6451.t233 a_5396_8177.t4 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1549 AVDD.t73 AVDD.t72 AVDD.t73 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1550 a_n13990_n5465.t114 a_n11737_n14973.t101 AVSS.t341 AVSS.t144 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1551 a_n13990_8177.t108 IREF.t251 AVDD.t1416 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1552 AVSS.t35 AVSS.t33 AVSS.t35 AVSS.t34 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1553 a_n13990_8177.t336 VN.t83 a_n13990_n5465.t29 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1554 a_n13990_8177.t107 IREF.t252 AVDD.t1417 AVDD.t98 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1555 a_n11737_n14973.t9 IREF.t253 AVDD.t1418 AVDD.t480 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1556 a_n13990_n5465.t115 a_n11737_n14973.t102 AVSS.t342 AVSS.t141 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1557 a_n13990_8177.t78 VN.t84 a_n13990_n5465.t28 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1558 a_5396_8177.t92 a_n11317_n20927.t1 a_5396_n6451.t7 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1559 AVDD.t71 AVDD.t69 AVDD.t71 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1560 AVDD.t68 AVDD.t66 AVDD.t68 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1561 AVDD.t1281 IREF.t0 IREF.t1 AVDD.t810 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1562 a_n13990_n6451.t54 VP.t87 a_n13990_8177.t62 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1563 a_n13990_n6451.t28 a_n11737_n14973.t103 AVSS.t343 AVSS.t82 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1564 AVDD.t1419 IREF.t254 a_n13990_8177.t106 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1565 AVSS.t32 AVSS.t30 AVSS.t32 AVSS.t31 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X1566 AVSS.t29 AVSS.t27 AVSS.t29 AVSS.t28 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1567 AVDD.t65 AVDD.t64 AVDD.t65 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1568 AVDD.t63 AVDD.t61 AVDD.t63 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1569 AVDD.t60 AVDD.t58 AVDD.t60 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1570 AVDD.t57 AVDD.t55 AVDD.t57 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1571 a_5396_9163.t4 a_5396_n6451.t234 AVDD.t1519 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1572 AVDD.t54 AVDD.t52 AVDD.t54 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1573 a_n13990_8177.t79 VN.t85 a_n13990_n5465.t27 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1574 a_5396_n6451.t43 a_n11317_n20927.t1 a_5396_8177.t91 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1575 AVDD.t1520 a_5396_n6451.t235 a_5396_9163.t3 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1576 a_n13990_8177.t105 IREF.t255 AVDD.t1420 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1577 AVDD.t51 AVDD.t50 AVDD.t51 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1578 a_n13990_8177.t104 IREF.t256 AVDD.t1421 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1579 a_5396_8177.t90 a_n11317_n20927.t1 a_5396_n6451.t20 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1580 AVDD.t49 AVDD.t48 AVDD.t49 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1581 AVSS.t26 AVSS.t24 AVSS.t26 AVSS.t25 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1582 VOUT.t2 a_n11317_n20927.t1 a_5396_9163.t118 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1583 a_n13990_n5465.t26 VN.t86 a_n13990_8177.t80 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1584 a_5396_9163.t2 a_5396_n6451.t236 AVDD.t1521 AVDD.t111 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1585 AVSS.t23 AVSS.t21 AVSS.t23 AVSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1586 a_5396_8177.t3 a_5396_n6451.t237 AVDD.t1522 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1587 AVSS.t20 AVSS.t18 AVSS.t20 AVSS.t19 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1588 AVSS.t17 AVSS.t15 AVSS.t17 AVSS.t16 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1589 AVSS.t14 AVSS.t12 AVSS.t14 AVSS.t13 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1590 AVDD.t47 AVDD.t46 AVDD.t47 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1591 AVSS.t11 AVSS.t9 AVSS.t11 AVSS.t10 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1592 AVDD.t45 AVDD.t43 AVDD.t45 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1593 a_n13990_8177.t103 IREF.t257 AVDD.t1422 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1594 a_n13990_8177.t102 IREF.t258 AVDD.t1423 AVDD.t205 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1595 VOUT.t1 a_n11317_n20927.t1 a_5396_9163.t163 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1596 AVDD.t42 AVDD.t41 AVDD.t42 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1597 AVDD.t40 AVDD.t38 AVDD.t40 AVDD.t39 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1598 AVDD.t37 AVDD.t35 AVDD.t37 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1599 AVDD.t34 AVDD.t32 AVDD.t34 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1600 a_5396_8177.t2 a_5396_n6451.t238 AVDD.t1523 AVDD.t193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1601 a_5396_8177.t89 a_n11317_n20927.t1 a_5396_n6451.t42 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1602 a_5396_9163.t1 a_5396_n6451.t239 AVDD.t1524 AVDD.t175 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1603 a_n13990_8177.t101 IREF.t259 AVDD.t1424 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1604 AVSS.t8 AVSS.t6 AVSS.t8 AVSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1605 AVDD.t1425 IREF.t260 a_n13990_8177.t100 AVDD.t186 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1606 a_n11737_n14973.t8 IREF.t261 AVDD.t1426 AVDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1607 AVSS.t5 AVSS.t3 AVSS.t5 AVSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1608 AVDD.t31 AVDD.t29 AVDD.t31 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1609 AVDD.t28 AVDD.t26 AVDD.t28 AVDD.t27 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1610 AVDD.t25 AVDD.t24 AVDD.t25 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1611 AVDD.t23 AVDD.t21 AVDD.t23 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1612 AVDD.t20 AVDD.t18 AVDD.t20 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1613 VOUT.t0 a_n11317_n20927.t1 a_5396_9163.t162 AVDD.t119 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1614 AVDD.t17 AVDD.t15 AVDD.t17 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1615 AVDD.t14 AVDD.t12 AVDD.t14 AVDD.t13 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1616 AVDD.t11 AVDD.t10 AVDD.t11 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1617 AVSS.t2 AVSS.t0 AVSS.t2 AVSS.t1 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1618 a_n13990_n5465.t5 a_n11737_n14973.t104 AVSS.t303 AVSS.t175 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1619 AVDD.t9 AVDD.t7 AVDD.t9 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1620 a_n13990_n5465.t25 VN.t87 a_n13990_8177.t81 AVDD.t93 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1621 a_5396_9163.t0 a_5396_n6451.t240 AVDD.t1525 AVDD.t178 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1622 a_n13990_n5465.t6 a_n11737_n14973.t105 AVSS.t304 AVSS.t172 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1623 AVDD.t6 AVDD.t4 AVDD.t6 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1624 a_n13990_8177.t99 IREF.t262 AVDD.t1374 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1625 AVDD.t1526 a_5396_n6451.t241 a_5396_8177.t1 AVDD.t88 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1626 a_n13990_8177.t98 IREF.t263 AVDD.t1375 AVDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1627 AVDD.t3 AVDD.t1 AVDD.t3 AVDD.t2 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1628 a_5396_n6451.t41 a_n11317_n20927.t1 a_5396_8177.t88 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1629 a_5396_8177.t0 a_5396_n6451.t242 AVDD.t1527 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
R0 AVDD.n1054 AVDD.n896 714.056
R1 AVDD.n1054 AVDD.n895 712.232
R2 AVDD.n1059 AVDD.n896 707.59
R3 AVDD.n1059 AVDD.n895 705.766
R4 AVDD.n1218 AVDD.n41 647.574
R5 AVDD.n1943 AVDD.n4 647.574
R6 AVDD.n1395 AVDD.n1 647.574
R7 AVDD.n85 AVDD.n84 647.574
R8 AVDD.n23 AVDD.n21 647.574
R9 AVDD.n1364 AVDD.n105 647.574
R10 AVDD.n92 AVDD.n86 647.574
R11 AVDD.n1220 AVDD.n655 647.574
R12 AVDD.n825 AVDD.n9 647.574
R13 AVDD.n111 AVDD.n11 647.574
R14 AVDD.n441 AVDD.n87 647.574
R15 AVDD.n1154 AVDD.n658 647.574
R16 AVDD.n1978 AVDD.n20 647.574
R17 AVDD.n112 AVDD.n14 647.574
R18 AVDD.n509 AVDD.n88 647.574
R19 AVDD.n656 AVDD.n36 647.574
R20 AVDD.n1950 AVDD.n41 642.269
R21 AVDD.n2017 AVDD.n4 642.269
R22 AVDD.n1408 AVDD.n1395 642.269
R23 AVDD.n85 AVDD.n83 642.269
R24 AVDD.n21 AVDD.n6 642.269
R25 AVDD.n1410 AVDD.n105 642.269
R26 AVDD.n91 AVDD.n86 642.269
R27 AVDD.n655 AVDD.n39 642.269
R28 AVDD.n2015 AVDD.n9 642.269
R29 AVDD.n111 AVDD.n108 642.269
R30 AVDD.n556 AVDD.n87 642.269
R31 AVDD.n658 AVDD.n38 642.269
R32 AVDD.n1978 AVDD.n7 642.269
R33 AVDD.n112 AVDD.n107 642.269
R34 AVDD.n554 AVDD.n88 642.269
R35 AVDD.n1952 AVDD.n36 642.269
R36 AVDD.n1218 AVDD.n40 640.197
R37 AVDD.n1943 AVDD.n3 640.197
R38 AVDD.n109 AVDD.n1 640.197
R39 AVDD.n1436 AVDD.n84 640.197
R40 AVDD.n1976 AVDD.n23 640.197
R41 AVDD.n1364 AVDD.n104 640.197
R42 AVDD.n1434 AVDD.n92 640.197
R43 AVDD.n1220 AVDD.n644 640.197
R44 AVDD.n825 AVDD.n8 640.197
R45 AVDD.n1393 AVDD.n11 640.197
R46 AVDD.n441 AVDD.n90 640.197
R47 AVDD.n1154 AVDD.n657 640.197
R48 AVDD.n22 AVDD.n20 640.197
R49 AVDD.n113 AVDD.n14 640.197
R50 AVDD.n509 AVDD.n89 640.197
R51 AVDD.n656 AVDD.n35 640.197
R52 AVDD.n1950 AVDD.n40 634.891
R53 AVDD.n2017 AVDD.n3 634.891
R54 AVDD.n1408 AVDD.n109 634.891
R55 AVDD.n1436 AVDD.n83 634.891
R56 AVDD.n1976 AVDD.n6 634.891
R57 AVDD.n1410 AVDD.n104 634.891
R58 AVDD.n1434 AVDD.n91 634.891
R59 AVDD.n644 AVDD.n39 634.891
R60 AVDD.n2015 AVDD.n8 634.891
R61 AVDD.n1393 AVDD.n108 634.891
R62 AVDD.n556 AVDD.n90 634.891
R63 AVDD.n657 AVDD.n38 634.891
R64 AVDD.n22 AVDD.n7 634.891
R65 AVDD.n113 AVDD.n107 634.891
R66 AVDD.n554 AVDD.n89 634.891
R67 AVDD.n1952 AVDD.n35 634.891
R68 AVDD.n979 AVDD.n898 351.805
R69 AVDD.n1052 AVDD.n898 351.639
R70 AVDD.n979 AVDD.n897 350.479
R71 AVDD.n1052 AVDD.n897 350.313
R72 AVDD.n355 AVDD.n140 322.38
R73 AVDD.n552 AVDD.n357 289.171
R74 AVDD.n316 AVDD.n141 289.171
R75 AVDD.n350 AVDD.n141 267.75
R76 AVDD.n357 AVDD.n355 255.06
R77 AVDD.n350 AVDD.n140 255.06
R78 AVDD.t328 AVDD.t13 85.1494
R79 AVDD.t131 AVDD.t39 85.1494
R80 AVDD.t810 AVDD.t181 85.1494
R81 AVDD.t373 AVDD.t2 81.7244
R82 AVDD.t638 AVDD.t875 79.7265
R83 AVDD.t2 AVDD.t264 79.5362
R84 AVDD.n1057 AVDD.t27 68.5002
R85 AVDD.t394 AVDD.t328 54.0391
R86 AVDD.t39 AVDD.t555 54.0391
R87 AVDD.t555 AVDD.t480 54.0391
R88 AVDD.t480 AVDD.t282 54.0391
R89 AVDD.t717 AVDD.t638 54.0391
R90 AVDD.t875 AVDD.t366 54.0391
R91 AVDD.t366 AVDD.t323 54.0391
R92 AVDD.t323 AVDD.t810 54.0391
R93 AVDD.t27 AVDD.n1055 50.3287
R94 AVDD.n2016 AVDD.n5 46.8594
R95 AVDD.n979 AVDD.t373 45.4522
R96 AVDD.t181 AVDD.n1054 45.3596
R97 AVDD.n1053 AVDD.t13 45.2864
R98 AVDD.n1058 AVDD.t131 45.2864
R99 AVDD.n978 AVDD.t394 37.9607
R100 AVDD.t67 AVDD.t44 31.8205
R101 AVDD.t79 AVDD.t241 31.8205
R102 AVDD.t178 AVDD.t56 31.8205
R103 AVDD.t22 AVDD.t114 31.8205
R104 AVDD.t294 AVDD.t70 31.8205
R105 AVDD.t16 AVDD.t335 31.8205
R106 AVDD.t33 AVDD.t62 31.8205
R107 AVDD.t347 AVDD.t381 29.7939
R108 AVDD.t193 AVDD.t59 29.7939
R109 AVDD.t200 AVDD.t226 29.7939
R110 AVDD.t156 AVDD.t338 29.7939
R111 AVDD.t5 AVDD.t153 29.7939
R112 AVDD.t0 AVDD.t252 29.7939
R113 AVDD.t82 AVDD.t238 29.7939
R114 AVDD.t233 AVDD.t93 29.7939
R115 AVDD.t44 AVDD.t19 20.1946
R116 AVDD.t19 AVDD.t122 20.1946
R117 AVDD.t122 AVDD.t347 20.1946
R118 AVDD.t59 AVDD.t88 20.1946
R119 AVDD.t279 AVDD.t193 20.1946
R120 AVDD.t291 AVDD.t279 20.1946
R121 AVDD.t241 AVDD.t291 20.1946
R122 AVDD.t148 AVDD.t178 20.1946
R123 AVDD.t111 AVDD.t148 20.1946
R124 AVDD.t226 AVDD.t111 20.1946
R125 AVDD.t175 AVDD.t156 20.1946
R126 AVDD.t338 AVDD.t399 20.1946
R127 AVDD.t399 AVDD.t119 20.1946
R128 AVDD.t119 AVDD.t22 20.1946
R129 AVDD.t141 AVDD.t294 20.1946
R130 AVDD.t136 AVDD.t141 20.1946
R131 AVDD.t153 AVDD.t136 20.1946
R132 AVDD.t252 AVDD.t98 20.1946
R133 AVDD.t53 AVDD.t0 20.1946
R134 AVDD.t30 AVDD.t53 20.1946
R135 AVDD.t335 AVDD.t30 20.1946
R136 AVDD.t205 AVDD.t255 20.1946
R137 AVDD.t255 AVDD.t36 20.1946
R138 AVDD.t36 AVDD.t82 20.1946
R139 AVDD.t186 AVDD.t233 20.1946
R140 AVDD.t93 AVDD.t378 20.1946
R141 AVDD.t378 AVDD.t85 20.1946
R142 AVDD.t85 AVDD.t33 20.1946
R143 AVDD.n1435 AVDD.t381 19.0569
R144 AVDD.n1394 AVDD.t200 19.0569
R145 AVDD.n1977 AVDD.t5 19.0569
R146 AVDD.t238 AVDD.n1056 19.0569
R147 AVDD.n555 AVDD.t67 16.9237
R148 AVDD.n106 AVDD.t79 16.9237
R149 AVDD.n1409 AVDD.t56 16.9237
R150 AVDD.t114 AVDD.n5 16.9237
R151 AVDD.n2016 AVDD.t70 16.9237
R152 AVDD.n37 AVDD.t16 16.9237
R153 AVDD.n1951 AVDD.t8 16.9237
R154 AVDD.n1219 AVDD.t62 16.9237
R155 AVDD.n1057 AVDD.t8 16.4971
R156 AVDD.t264 AVDD.n978 16.0789
R157 AVDD.n1057 AVDD.t205 15.3239
R158 AVDD.n1058 AVDD.n1053 13.7004
R159 AVDD.t282 AVDD.n1057 11.2268
R160 AVDD.n0 AVDD.t431 8.10567
R161 AVDD.n2021 AVDD.t953 8.10567
R162 AVDD.n2020 AVDD.t854 8.10567
R163 AVDD.n1352 AVDD.t923 8.10567
R164 AVDD.n1353 AVDD.t1105 8.10567
R165 AVDD.n1355 AVDD.t349 8.10567
R166 AVDD.n0 AVDD.t1187 8.10567
R167 AVDD.n2021 AVDD.t415 8.10567
R168 AVDD.n2020 AVDD.t320 8.10567
R169 AVDD.n1352 AVDD.t391 8.10567
R170 AVDD.n1353 AVDD.t587 8.10567
R171 AVDD.n1355 AVDD.t1083 8.10567
R172 AVDD.n1359 AVDD.t981 8.10567
R173 AVDD.n1361 AVDD.t207 8.10567
R174 AVDD.n1362 AVDD.t69 8.10567
R175 AVDD.n1367 AVDD.t211 8.10567
R176 AVDD.n1368 AVDD.t72 8.10567
R177 AVDD.n1370 AVDD.t676 8.10567
R178 AVDD.n1359 AVDD.t441 8.10567
R179 AVDD.n1361 AVDD.t959 8.10567
R180 AVDD.n1362 AVDD.t866 8.10567
R181 AVDD.n1367 AVDD.t221 8.10567
R182 AVDD.n1368 AVDD.t113 8.10567
R183 AVDD.n1370 AVDD.t694 8.10567
R184 AVDD.n1375 AVDD.t680 8.10567
R185 AVDD.n1373 AVDD.t1177 8.10567
R186 AVDD.n1372 AVDD.t1059 8.10567
R187 AVDD.n2012 AVDD.t1065 8.10567
R188 AVDD.n2011 AVDD.t759 8.10567
R189 AVDD.n2009 AVDD.t848 8.10567
R190 AVDD.n1375 AVDD.t702 8.10567
R191 AVDD.n1373 AVDD.t1191 8.10567
R192 AVDD.n1372 AVDD.t1069 8.10567
R193 AVDD.n2012 AVDD.t1089 8.10567
R194 AVDD.n2011 AVDD.t261 8.10567
R195 AVDD.n2009 AVDD.t314 8.10567
R196 AVDD.n2005 AVDD.t1225 8.10567
R197 AVDD.n2003 AVDD.t668 8.10567
R198 AVDD.n2002 AVDD.t793 8.10567
R199 AVDD.n1998 AVDD.t781 8.10567
R200 AVDD.n1997 AVDD.t889 8.10567
R201 AVDD.n1995 AVDD.t370 8.10567
R202 AVDD.n2005 AVDD.t725 8.10567
R203 AVDD.n2003 AVDD.t128 8.10567
R204 AVDD.n2002 AVDD.t266 8.10567
R205 AVDD.n1998 AVDD.t247 8.10567
R206 AVDD.n1997 AVDD.t353 8.10567
R207 AVDD.n1995 AVDD.t1119 8.10567
R208 AVDD.n68 AVDD.t138 8.10567
R209 AVDD.n67 AVDD.t1007 8.10567
R210 AVDD.n155 AVDD.t1263 8.10567
R211 AVDD.n152 AVDD.t421 8.10567
R212 AVDD.n151 AVDD.t383 8.10567
R213 AVDD.n162 AVDD.t670 8.10567
R214 AVDD.n150 AVDD.t1075 8.10567
R215 AVDD.n149 AVDD.t1107 8.10567
R216 AVDD.n170 AVDD.t110 8.10567
R217 AVDD.n147 AVDD.t652 8.10567
R218 AVDD.n146 AVDD.t933 8.10567
R219 AVDD.n45 AVDD.t1207 8.10567
R220 AVDD.n44 AVDD.t947 8.10567
R221 AVDD.n1614 AVDD.t52 8.10567
R222 AVDD.n1611 AVDD.t1063 8.10567
R223 AVDD.n1610 AVDD.t1135 8.10567
R224 AVDD.n1621 AVDD.t712 8.10567
R225 AVDD.n1609 AVDD.t417 8.10567
R226 AVDD.n1608 AVDD.t286 8.10567
R227 AVDD.n1629 AVDD.t268 8.10567
R228 AVDD.n65 AVDD.t642 8.10567
R229 AVDD.n64 AVDD.t1167 8.10567
R230 AVDD.n1938 AVDD.t46 8.10567
R231 AVDD.n1940 AVDD.t583 8.10567
R232 AVDD.n1941 AVDD.t451 8.10567
R233 AVDD.n1947 AVDD.t550 8.10567
R234 AVDD.n1946 AVDD.t751 8.10567
R235 AVDD.n1944 AVDD.t1235 8.10567
R236 AVDD.n1938 AVDD.t168 8.10567
R237 AVDD.n1940 AVDD.t690 8.10567
R238 AVDD.n1941 AVDD.t577 8.10567
R239 AVDD.n1947 AVDD.t650 8.10567
R240 AVDD.n1946 AVDD.t862 8.10567
R241 AVDD.n1944 AVDD.t48 8.10567
R242 AVDD.n1958 AVDD.t605 8.10567
R243 AVDD.n1956 AVDD.t1099 8.10567
R244 AVDD.n1955 AVDD.t999 8.10567
R245 AVDD.n1259 AVDD.t881 8.10567
R246 AVDD.n1260 AVDD.t773 8.10567
R247 AVDD.n1958 AVDD.t719 8.10567
R248 AVDD.n1956 AVDD.t1205 8.10567
R249 AVDD.n1955 AVDD.t1095 8.10567
R250 AVDD.n1259 AVDD.t457 8.10567
R251 AVDD.n1260 AVDD.t357 8.10567
R252 AVDD.n652 AVDD.t104 8.10567
R253 AVDD.n1230 AVDD.t664 8.10567
R254 AVDD.n650 AVDD.t284 8.10567
R255 AVDD.n1235 AVDD.t965 8.10567
R256 AVDD.n647 AVDD.t903 8.10567
R257 AVDD.n646 AVDD.t526 8.10567
R258 AVDD.n1242 AVDD.t905 8.10567
R259 AVDD.n642 AVDD.t500 8.10567
R260 AVDD.n1248 AVDD.t90 8.10567
R261 AVDD.n640 AVDD.t471 8.10567
R262 AVDD.n1253 AVDD.t747 8.10567
R263 AVDD.n637 AVDD.t1097 8.10567
R264 AVDD.n636 AVDD.t7 8.10567
R265 AVDD.n634 AVDD.t937 8.10567
R266 AVDD.n1266 AVDD.t1157 8.10567
R267 AVDD.n632 AVDD.t1067 8.10567
R268 AVDD.n1271 AVDD.t494 8.10567
R269 AVDD.n629 AVDD.t425 8.10567
R270 AVDD.n628 AVDD.t1015 8.10567
R271 AVDD.n1278 AVDD.t97 8.10567
R272 AVDD.n625 AVDD.t4 8.10567
R273 AVDD.n1284 AVDD.t593 8.10567
R274 AVDD.n623 AVDD.t1035 8.10567
R275 AVDD.n1289 AVDD.t1125 8.10567
R276 AVDD.n620 AVDD.t1209 8.10567
R277 AVDD.n652 AVDD.t116 8.10567
R278 AVDD.n1230 AVDD.t672 8.10567
R279 AVDD.n650 AVDD.t288 8.10567
R280 AVDD.n1235 AVDD.t971 8.10567
R281 AVDD.n647 AVDD.t909 8.10567
R282 AVDD.n646 AVDD.t532 8.10567
R283 AVDD.n1242 AVDD.t911 8.10567
R284 AVDD.n642 AVDD.t508 8.10567
R285 AVDD.n1248 AVDD.t102 8.10567
R286 AVDD.n640 AVDD.t484 8.10567
R287 AVDD.n1253 AVDD.t755 8.10567
R288 AVDD.n637 AVDD.t1103 8.10567
R289 AVDD.n636 AVDD.t24 8.10567
R290 AVDD.n634 AVDD.t941 8.10567
R291 AVDD.n1266 AVDD.t1165 8.10567
R292 AVDD.n632 AVDD.t1081 8.10567
R293 AVDD.n1271 AVDD.t502 8.10567
R294 AVDD.n629 AVDD.t429 8.10567
R295 AVDD.n628 AVDD.t1019 8.10567
R296 AVDD.n1278 AVDD.t106 8.10567
R297 AVDD.n625 AVDD.t10 8.10567
R298 AVDD.n1284 AVDD.t599 8.10567
R299 AVDD.n623 AVDD.t1045 8.10567
R300 AVDD.n1289 AVDD.t1133 8.10567
R301 AVDD.n620 AVDD.t1215 8.10567
R302 AVDD.n1224 AVDD.t625 8.10567
R303 AVDD.n1223 AVDD.t514 8.10567
R304 AVDD.n747 AVDD.t520 8.10567
R305 AVDD.n748 AVDD.t1195 8.10567
R306 AVDD.n1210 AVDD.t1129 8.10567
R307 AVDD.n1209 AVDD.t1013 8.10567
R308 AVDD.n1205 AVDD.t935 8.10567
R309 AVDD.n1204 AVDD.t832 8.10567
R310 AVDD.n1160 AVDD.t1245 8.10567
R311 AVDD.n1161 AVDD.t714 8.10567
R312 AVDD.n1162 AVDD.t765 8.10567
R313 AVDD.n1163 AVDD.t1169 8.10567
R314 AVDD.n1164 AVDD.t899 8.10567
R315 AVDD.n1165 AVDD.t619 8.10567
R316 AVDD.n1166 AVDD.t185 8.10567
R317 AVDD.n1167 AVDD.t237 8.10567
R318 AVDD.n1169 AVDD.t488 8.10567
R319 AVDD.n1170 AVDD.t35 8.10567
R320 AVDD.n1171 AVDD.t627 8.10567
R321 AVDD.n1172 AVDD.t204 8.10567
R322 AVDD.n1155 AVDD.t61 8.10567
R323 AVDD.n1157 AVDD.t595 8.10567
R324 AVDD.n1158 AVDD.t486 8.10567
R325 AVDD.n1215 AVDD.t563 8.10567
R326 AVDD.n1214 AVDD.t775 8.10567
R327 AVDD.n55 AVDD.t818 8.10567
R328 AVDD.n1779 AVDD.t868 8.10567
R329 AVDD.n57 AVDD.t1247 8.10567
R330 AVDD.n1774 AVDD.t995 8.10567
R331 AVDD.n58 AVDD.t731 8.10567
R332 AVDD.n1769 AVDD.t304 8.10567
R333 AVDD.n59 AVDD.t342 8.10567
R334 AVDD.n60 AVDD.t585 8.10567
R335 AVDD.n1761 AVDD.t145 8.10567
R336 AVDD.n61 AVDD.t737 8.10567
R337 AVDD.n62 AVDD.t310 8.10567
R338 AVDD.n1962 AVDD.t1111 8.10567
R339 AVDD.n30 AVDD.t852 8.10567
R340 AVDD.n1967 AVDD.t1241 8.10567
R341 AVDD.n27 AVDD.t987 8.10567
R342 AVDD.n26 AVDD.t1023 8.10567
R343 AVDD.n1974 AVDD.t609 8.10567
R344 AVDD.n1299 AVDD.t330 8.10567
R345 AVDD.n1303 AVDD.t152 8.10567
R346 AVDD.n1296 AVDD.t135 8.10567
R347 AVDD.n1308 AVDD.t548 8.10567
R348 AVDD.n1293 AVDD.t1055 8.10567
R349 AVDD.n1962 AVDD.t465 8.10567
R350 AVDD.n30 AVDD.t188 8.10567
R351 AVDD.n1967 AVDD.t617 8.10567
R352 AVDD.n27 AVDD.t340 8.10567
R353 AVDD.n26 AVDD.t375 8.10567
R354 AVDD.n1974 AVDD.t1227 8.10567
R355 AVDD.n1299 AVDD.t963 8.10567
R356 AVDD.n1303 AVDD.t812 8.10567
R357 AVDD.n1296 AVDD.t799 8.10567
R358 AVDD.n1308 AVDD.t1173 8.10567
R359 AVDD.n1293 AVDD.t411 8.10567
R360 AVDD.n449 AVDD.t735 8.10567
R361 AVDD.n450 AVDD.t1163 8.10567
R362 AVDD.n451 AVDD.t278 8.10567
R363 AVDD.n452 AVDD.t698 8.10567
R364 AVDD.n453 AVDD.t969 8.10567
R365 AVDD.n454 AVDD.t1233 8.10567
R366 AVDD.n455 AVDD.t380 8.10567
R367 AVDD.n457 AVDD.t346 8.10567
R368 AVDD.n458 AVDD.t623 8.10567
R369 AVDD.n459 AVDD.t939 8.10567
R370 AVDD.n460 AVDD.t1199 8.10567
R371 AVDD.n461 AVDD.t150 8.10567
R372 AVDD.n449 AVDD.t1139 8.10567
R373 AVDD.n450 AVDD.t290 8.10567
R374 AVDD.n451 AVDD.t674 8.10567
R375 AVDD.n452 AVDD.t1077 8.10567
R376 AVDD.n453 AVDD.t58 8.10567
R377 AVDD.n454 AVDD.t363 8.10567
R378 AVDD.n455 AVDD.t803 8.10567
R379 AVDD.n457 AVDD.t757 8.10567
R380 AVDD.n458 AVDD.t1021 8.10567
R381 AVDD.n459 AVDD.t18 8.10567
R382 AVDD.n460 AVDD.t332 8.10567
R383 AVDD.n461 AVDD.t569 8.10567
R384 AVDD.n411 AVDD.t557 8.10567
R385 AVDD.n409 AVDD.t118 8.10567
R386 AVDD.n416 AVDD.t398 8.10567
R387 AVDD.n406 AVDD.t838 8.10567
R388 AVDD.n405 AVDD.t795 8.10567
R389 AVDD.n423 AVDD.t1051 8.10567
R390 AVDD.n402 AVDD.t199 8.10567
R391 AVDD.n429 AVDD.t225 8.10567
R392 AVDD.n400 AVDD.t504 8.10567
R393 AVDD.n434 AVDD.t1029 8.10567
R394 AVDD.n397 AVDD.t1279 8.10567
R395 AVDD.n411 AVDD.t949 8.10567
R396 AVDD.n409 AVDD.t522 8.10567
R397 AVDD.n416 AVDD.t814 8.10567
R398 AVDD.n406 AVDD.t1217 8.10567
R399 AVDD.n405 AVDD.t1175 8.10567
R400 AVDD.n423 AVDD.t174 8.10567
R401 AVDD.n402 AVDD.t611 8.10567
R402 AVDD.n429 AVDD.t629 8.10567
R403 AVDD.n400 AVDD.t915 8.10567
R404 AVDD.n434 AVDD.t147 8.10567
R405 AVDD.n397 AVDD.t433 8.10567
R406 AVDD.n467 AVDD.t1255 8.10567
R407 AVDD.n466 AVDD.t100 8.10567
R408 AVDD.n550 AVDD.t66 8.10567
R409 AVDD.n549 AVDD.t202 8.10567
R410 AVDD.n547 AVDD.t979 8.10567
R411 AVDD.n560 AVDD.t1093 8.10567
R412 AVDD.n559 AVDD.t997 8.10567
R413 AVDD.n463 AVDD.t1003 8.10567
R414 AVDD.n464 AVDD.t635 8.10567
R415 AVDD.n1379 AVDD.t453 8.10567
R416 AVDD.n618 AVDD.t1039 8.10567
R417 AVDD.n1384 AVDD.t1109 8.10567
R418 AVDD.n615 AVDD.t761 8.10567
R419 AVDD.n116 AVDD.t155 8.10567
R420 AVDD.n1391 AVDD.t230 8.10567
R421 AVDD.n612 AVDD.t1145 8.10567
R422 AVDD.n117 AVDD.t461 8.10567
R423 AVDD.n118 AVDD.t534 8.10567
R424 AVDD.n119 AVDD.t164 8.10567
R425 AVDD.n120 AVDD.t243 8.10567
R426 AVDD.n121 AVDD.t967 8.10567
R427 AVDD.n126 AVDD.t407 8.10567
R428 AVDD.n127 AVDD.t1147 8.10567
R429 AVDD.n128 AVDD.t785 8.10567
R430 AVDD.n129 AVDD.t856 8.10567
R431 AVDD.n130 AVDD.t459 8.10567
R432 AVDD.n131 AVDD.t858 8.10567
R433 AVDD.n132 AVDD.t907 8.10567
R434 AVDD.n133 AVDD.t530 8.10567
R435 AVDD.n135 AVDD.t1223 8.10567
R436 AVDD.n136 AVDD.t1269 8.10567
R437 AVDD.n137 AVDD.t767 8.10567
R438 AVDD.n138 AVDD.t820 8.10567
R439 AVDD.n139 AVDD.t591 8.10567
R440 AVDD.n1379 AVDD.t463 8.10567
R441 AVDD.n618 AVDD.t1047 8.10567
R442 AVDD.n1384 AVDD.t1117 8.10567
R443 AVDD.n615 AVDD.t769 8.10567
R444 AVDD.n116 AVDD.t160 8.10567
R445 AVDD.n1391 AVDD.t235 8.10567
R446 AVDD.n612 AVDD.t1151 8.10567
R447 AVDD.n117 AVDD.t473 8.10567
R448 AVDD.n118 AVDD.t540 8.10567
R449 AVDD.n119 AVDD.t172 8.10567
R450 AVDD.n120 AVDD.t249 8.10567
R451 AVDD.n121 AVDD.t975 8.10567
R452 AVDD.n126 AVDD.t409 8.10567
R453 AVDD.n127 AVDD.t1155 8.10567
R454 AVDD.n128 AVDD.t787 8.10567
R455 AVDD.n129 AVDD.t864 8.10567
R456 AVDD.n130 AVDD.t467 8.10567
R457 AVDD.n131 AVDD.t860 8.10567
R458 AVDD.n132 AVDD.t913 8.10567
R459 AVDD.n133 AVDD.t538 8.10567
R460 AVDD.n135 AVDD.t1229 8.10567
R461 AVDD.n136 AVDD.t1273 8.10567
R462 AVDD.n137 AVDD.t771 8.10567
R463 AVDD.n138 AVDD.t828 8.10567
R464 AVDD.n139 AVDD.t597 8.10567
R465 AVDD.n438 AVDD.t197 8.10567
R466 AVDD.n439 AVDD.t55 8.10567
R467 AVDD.n444 AVDD.t74 8.10567
R468 AVDD.n445 AVDD.t546 8.10567
R469 AVDD.n447 AVDD.t603 8.10567
R470 AVDD.n438 AVDD.t929 8.10567
R471 AVDD.n439 AVDD.t824 8.10567
R472 AVDD.n444 AVDD.t842 8.10567
R473 AVDD.n445 AVDD.t830 8.10567
R474 AVDD.n447 AVDD.t162 8.10567
R475 AVDD.n504 AVDD.t1001 8.10567
R476 AVDD.n506 AVDD.t419 8.10567
R477 AVDD.n507 AVDD.t544 8.10567
R478 AVDD.n512 AVDD.t528 8.10567
R479 AVDD.n513 AVDD.t633 8.10567
R480 AVDD.n515 AVDD.t126 8.10567
R481 AVDD.n504 AVDD.t581 8.10567
R482 AVDD.n506 AVDD.t1257 8.10567
R483 AVDD.n507 AVDD.t108 8.10567
R484 AVDD.n512 AVDD.t78 8.10567
R485 AVDD.n513 AVDD.t213 8.10567
R486 AVDD.n515 AVDD.t989 8.10567
R487 AVDD.n519 AVDD.t274 8.10567
R488 AVDD.n363 AVDD.t688 8.10567
R489 AVDD.n524 AVDD.t1061 8.10567
R490 AVDD.n362 AVDD.t217 8.10567
R491 AVDD.n361 AVDD.t490 8.10567
R492 AVDD.n531 AVDD.t791 8.10567
R493 AVDD.n360 AVDD.t1189 8.10567
R494 AVDD.n537 AVDD.t1159 8.10567
R495 AVDD.n359 AVDD.t133 8.10567
R496 AVDD.n542 AVDD.t445 8.10567
R497 AVDD.n358 AVDD.t749 8.10567
R498 AVDD.n370 AVDD.t50 8.10567
R499 AVDD.n369 AVDD.t943 8.10567
R500 AVDD.n375 AVDD.t1201 8.10567
R501 AVDD.n368 AVDD.t359 8.10567
R502 AVDD.n367 AVDD.t316 8.10567
R503 AVDD.n382 AVDD.t589 8.10567
R504 AVDD.n366 AVDD.t1011 8.10567
R505 AVDD.n388 AVDD.t1027 8.10567
R506 AVDD.n365 AVDD.t1277 8.10567
R507 AVDD.n393 AVDD.t579 8.10567
R508 AVDD.n364 AVDD.t872 8.10567
R509 AVDD.n1397 AVDD.t209 8.10567
R510 AVDD.n1399 AVDD.t729 8.10567
R511 AVDD.n1400 AVDD.t607 8.10567
R512 AVDD.n1405 AVDD.t684 8.10567
R513 AVDD.n1404 AVDD.t893 8.10567
R514 AVDD.n1402 AVDD.t95 8.10567
R515 AVDD.n1397 AVDD.t1049 8.10567
R516 AVDD.n1399 AVDD.t300 8.10567
R517 AVDD.n1400 AVDD.t166 8.10567
R518 AVDD.n1405 AVDD.t270 8.10567
R519 AVDD.n1404 AVDD.t439 8.10567
R520 AVDD.n1402 AVDD.t957 8.10567
R521 AVDD.n1416 AVDD.t753 8.10567
R522 AVDD.n1414 AVDD.t1237 8.10567
R523 AVDD.n1413 AVDD.t1143 8.10567
R524 AVDD.n122 AVDD.t498 8.10567
R525 AVDD.n123 AVDD.t389 8.10567
R526 AVDD.n1416 AVDD.t318 8.10567
R527 AVDD.n1414 AVDD.t836 8.10567
R528 AVDD.n1413 AVDD.t721 8.10567
R529 AVDD.n122 AVDD.t1219 8.10567
R530 AVDD.n123 AVDD.t1115 8.10567
R531 AVDD.n1420 AVDD.t240 8.10567
R532 AVDD.n99 AVDD.t660 8.10567
R533 AVDD.n1425 AVDD.t1033 8.10567
R534 AVDD.n96 AVDD.t192 8.10567
R535 AVDD.n95 AVDD.t455 8.10567
R536 AVDD.n1432 AVDD.t763 8.10567
R537 AVDD.n329 AVDD.t1171 8.10567
R538 AVDD.n333 AVDD.t1127 8.10567
R539 AVDD.n326 AVDD.t121 8.10567
R540 AVDD.n338 AVDD.t423 8.10567
R541 AVDD.n323 AVDD.t727 8.10567
R542 AVDD.n343 AVDD.t951 8.10567
R543 AVDD.n1420 AVDD.t885 8.10567
R544 AVDD.n99 AVDD.t1267 8.10567
R545 AVDD.n1425 AVDD.t403 8.10567
R546 AVDD.n96 AVDD.t846 8.10567
R547 AVDD.n95 AVDD.t1091 8.10567
R548 AVDD.n1432 AVDD.t87 8.10567
R549 AVDD.n329 AVDD.t524 8.10567
R550 AVDD.n333 AVDD.t482 8.10567
R551 AVDD.n326 AVDD.t777 8.10567
R552 AVDD.n338 AVDD.t1057 8.10567
R553 AVDD.n323 AVDD.t43 8.10567
R554 AVDD.n343 AVDD.t308 8.10567
R555 AVDD.n346 AVDD.t822 8.10567
R556 AVDD.n347 AVDD.t710 8.10567
R557 AVDD.n352 AVDD.t124 8.10567
R558 AVDD.n353 AVDD.t1271 8.10567
R559 AVDD.n311 AVDD.t1037 8.10567
R560 AVDD.n313 AVDD.t296 8.10567
R561 AVDD.n314 AVDD.t158 8.10567
R562 AVDD.n319 AVDD.t259 8.10567
R563 AVDD.n320 AVDD.t427 8.10567
R564 AVDD.n78 AVDD.t344 8.10567
R565 AVDD.n1448 AVDD.t779 8.10567
R566 AVDD.n80 AVDD.t1161 8.10567
R567 AVDD.n1443 AVDD.t306 8.10567
R568 AVDD.n81 AVDD.t575 8.10567
R569 AVDD.n1438 AVDD.t870 8.10567
R570 AVDD.n297 AVDD.t1253 8.10567
R571 AVDD.n301 AVDD.t1213 8.10567
R572 AVDD.n296 AVDD.t223 8.10567
R573 AVDD.n306 AVDD.t536 8.10567
R574 AVDD.n142 AVDD.t826 8.10567
R575 AVDD.n1312 AVDD.t21 8.10567
R576 AVDD.n1313 AVDD.t917 8.10567
R577 AVDD.n1314 AVDD.t1181 8.10567
R578 AVDD.n1315 AVDD.t337 8.10567
R579 AVDD.n1316 AVDD.t298 8.10567
R580 AVDD.n1317 AVDD.t567 8.10567
R581 AVDD.n1318 AVDD.t993 8.10567
R582 AVDD.n1319 AVDD.t1009 8.10567
R583 AVDD.n1320 AVDD.t1265 8.10567
R584 AVDD.n1321 AVDD.t559 8.10567
R585 AVDD.n1322 AVDD.t844 8.10567
R586 AVDD.n1312 AVDD.t692 8.10567
R587 AVDD.n1313 AVDD.t276 8.10567
R588 AVDD.n1314 AVDD.t552 8.10567
R589 AVDD.n1315 AVDD.t973 8.10567
R590 AVDD.n1316 AVDD.t927 8.10567
R591 AVDD.n1317 AVDD.t1193 8.10567
R592 AVDD.n1318 AVDD.t351 8.10567
R593 AVDD.n1319 AVDD.t368 8.10567
R594 AVDD.n1320 AVDD.t648 8.10567
R595 AVDD.n1321 AVDD.t1179 8.10567
R596 AVDD.n1322 AVDD.t177 8.10567
R597 AVDD.n959 AVDD.t1079 8.10567
R598 AVDD.n936 AVDD.t658 8.10567
R599 AVDD.n899 AVDD.t783 8.10567
R600 AVDD.n926 AVDD.t190 8.10567
R601 AVDD.n1121 AVDD.t945 8.10567
R602 AVDD.n1120 AVDD.t130 8.10567
R603 AVDD.n665 AVDD.t678 8.10567
R604 AVDD.n1136 AVDD.t1185 8.10567
R605 AVDD.n711 AVDD.t921 8.10567
R606 AVDD.n715 AVDD.t640 8.10567
R607 AVDD.n705 AVDD.t215 8.10567
R608 AVDD.n700 AVDD.t272 8.10567
R609 AVDD.n888 AVDD.t510 8.10567
R610 AVDD.n697 AVDD.t64 8.10567
R611 AVDD.n725 AVDD.t656 8.10567
R612 AVDD.n724 AVDD.t228 8.10567
R613 AVDD.n728 AVDD.t1249 8.10567
R614 AVDD.n846 AVDD.t76 8.10567
R615 AVDD.n862 AVDD.t1153 8.10567
R616 AVDD.n859 AVDD.t879 8.10567
R617 AVDD.n1138 AVDD.t654 8.10567
R618 AVDD.n709 AVDD.t1203 8.10567
R619 AVDD.n716 AVDD.t743 8.10567
R620 AVDD.n701 AVDD.t365 8.10567
R621 AVDD.n702 AVDD.t1251 8.10567
R622 AVDD.n889 AVDD.t1043 8.10567
R623 AVDD.n696 AVDD.t1121 8.10567
R624 AVDD.n726 AVDD.t26 8.10567
R625 AVDD.n727 AVDD.t686 8.10567
R626 AVDD.n875 AVDD.t901 8.10567
R627 AVDD.n847 AVDD.t961 8.10567
R628 AVDD.n868 AVDD.t475 8.10567
R629 AVDD.n863 AVDD.t615 8.10567
R630 AVDD.n660 AVDD.t739 8.10567
R631 AVDD.n1143 AVDD.t789 8.10567
R632 AVDD.n745 AVDD.t312 8.10567
R633 AVDD.n744 AVDD.t413 8.10567
R634 AVDD.n1151 AVDD.t405 8.10567
R635 AVDD.n1150 AVDD.t516 8.10567
R636 AVDD.n1148 AVDD.t1261 8.10567
R637 AVDD.n857 AVDD.t1259 8.10567
R638 AVDD.n849 AVDD.t1005 8.10567
R639 AVDD.n850 AVDD.t1041 8.10567
R640 AVDD.n19 AVDD.t631 8.10567
R641 AVDD.n18 AVDD.t355 8.10567
R642 AVDD.n1984 AVDD.t183 8.10567
R643 AVDD.n17 AVDD.t170 8.10567
R644 AVDD.n1989 AVDD.t571 8.10567
R645 AVDD.n16 AVDD.t1073 8.10567
R646 AVDD.n822 AVDD.t565 8.10567
R647 AVDD.n823 AVDD.t437 8.10567
R648 AVDD.n828 AVDD.t449 8.10567
R649 AVDD.n829 AVDD.t1017 8.10567
R650 AVDD.n831 AVDD.t447 8.10567
R651 AVDD.n822 AVDD.t143 8.10567
R652 AVDD.n823 AVDD.t15 8.10567
R653 AVDD.n828 AVDD.t41 8.10567
R654 AVDD.n829 AVDD.t700 8.10567
R655 AVDD.n831 AVDD.t573 8.10567
R656 AVDD.n835 AVDD.t877 8.10567
R657 AVDD.n837 AVDD.t302 8.10567
R658 AVDD.n838 AVDD.t401 8.10567
R659 AVDD.n842 AVDD.t385 8.10567
R660 AVDD.n843 AVDD.t496 8.10567
R661 AVDD.n835 AVDD.t977 8.10567
R662 AVDD.n837 AVDD.t396 8.10567
R663 AVDD.n838 AVDD.t512 8.10567
R664 AVDD.n842 AVDD.t492 8.10567
R665 AVDD.n843 AVDD.t613 8.10567
R666 AVDD.n781 AVDD.t334 8.10567
R667 AVDD.n782 AVDD.t29 8.10567
R668 AVDD.n783 AVDD.t469 8.10567
R669 AVDD.n784 AVDD.t195 8.10567
R670 AVDD.n785 AVDD.t251 8.10567
R671 AVDD.n786 AVDD.t1085 8.10567
R672 AVDD.n787 AVDD.t834 8.10567
R673 AVDD.n789 AVDD.t662 8.10567
R674 AVDD.n790 AVDD.t644 8.10567
R675 AVDD.n791 AVDD.t1025 8.10567
R676 AVDD.n792 AVDD.t293 8.10567
R677 AVDD.n781 AVDD.t745 8.10567
R678 AVDD.n782 AVDD.t443 8.10567
R679 AVDD.n783 AVDD.t891 8.10567
R680 AVDD.n784 AVDD.t601 8.10567
R681 AVDD.n785 AVDD.t646 8.10567
R682 AVDD.n786 AVDD.t219 8.10567
R683 AVDD.n787 AVDD.t1211 8.10567
R684 AVDD.n789 AVDD.t1053 8.10567
R685 AVDD.n790 AVDD.t1031 8.10567
R686 AVDD.n791 AVDD.t140 8.10567
R687 AVDD.n792 AVDD.t682 8.10567
R688 AVDD.n743 AVDD.t477 8.10567
R689 AVDD.n754 AVDD.t1197 8.10567
R690 AVDD.n741 AVDD.t1231 8.10567
R691 AVDD.n759 AVDD.t377 8.10567
R692 AVDD.n738 AVDD.t92 8.10567
R693 AVDD.n737 AVDD.t1101 8.10567
R694 AVDD.n766 AVDD.t696 8.10567
R695 AVDD.n734 AVDD.t733 8.10567
R696 AVDD.n772 AVDD.t985 8.10567
R697 AVDD.n732 AVDD.t561 8.10567
R698 AVDD.n777 AVDD.t1123 8.10567
R699 AVDD.n729 AVDD.t708 8.10567
R700 AVDD.n743 AVDD.t895 8.10567
R701 AVDD.n754 AVDD.t325 8.10567
R702 AVDD.n741 AVDD.t361 8.10567
R703 AVDD.n759 AVDD.t801 8.10567
R704 AVDD.n738 AVDD.t506 8.10567
R705 AVDD.n737 AVDD.t232 8.10567
R706 AVDD.n766 AVDD.t1071 8.10567
R707 AVDD.n734 AVDD.t1137 8.10567
R708 AVDD.n772 AVDD.t81 8.10567
R709 AVDD.n732 AVDD.t955 8.10567
R710 AVDD.n777 AVDD.t254 8.10567
R711 AVDD.n729 AVDD.t1087 8.10567
R712 AVDD.n683 AVDD.t983 8.10567
R713 AVDD.n684 AVDD.t180 8.10567
R714 AVDD.n1098 AVDD.t723 8.10567
R715 AVDD.n942 AVDD.t1141 8.10567
R716 AVDD.n944 AVDD.t706 8.10567
R717 AVDD.n943 AVDD.t816 8.10567
R718 AVDD.n1027 AVDD.t245 8.10567
R719 AVDD.n919 AVDD.t809 8.10567
R720 AVDD.n1022 AVDD.t322 8.10567
R721 AVDD.n920 AVDD.t1221 8.10567
R722 AVDD.n1017 AVDD.t874 8.10567
R723 AVDD.n921 AVDD.t637 8.10567
R724 AVDD.n1012 AVDD.t716 8.10567
R725 AVDD.n922 AVDD.t925 8.10567
R726 AVDD.n923 AVDD.t281 8.10567
R727 AVDD.n1004 AVDD.t479 8.10567
R728 AVDD.n924 AVDD.t554 8.10567
R729 AVDD.n999 AVDD.t38 8.10567
R730 AVDD.n1160 AVDD.t621 8.10567
R731 AVDD.n1161 AVDD.t32 8.10567
R732 AVDD.n1162 AVDD.t84 8.10567
R733 AVDD.n1163 AVDD.t518 8.10567
R734 AVDD.n1164 AVDD.t257 8.10567
R735 AVDD.n1165 AVDD.t1239 8.10567
R736 AVDD.n1166 AVDD.t840 8.10567
R737 AVDD.n1167 AVDD.t883 8.10567
R738 AVDD.n1169 AVDD.t1113 8.10567
R739 AVDD.n1170 AVDD.t704 8.10567
R740 AVDD.n1171 AVDD.t1243 8.10567
R741 AVDD.n1172 AVDD.t850 8.10567
R742 AVDD.n934 AVDD.t327 6.64567
R743 AVDD.n966 AVDD.t393 6.64567
R744 AVDD.n932 AVDD.t1183 6.64567
R745 AVDD.n931 AVDD.t991 6.64567
R746 AVDD.n973 AVDD.t1275 6.64567
R747 AVDD.n975 AVDD.t919 6.64567
R748 AVDD.n976 AVDD.t542 6.64567
R749 AVDD.n976 AVDD.t887 6.64567
R750 AVDD.n982 AVDD.t807 6.64567
R751 AVDD.n982 AVDD.t1131 6.64567
R752 AVDD.n983 AVDD.t435 6.64567
R753 AVDD.n983 AVDD.t797 6.64567
R754 AVDD.n985 AVDD.t1 6.64567
R755 AVDD.n985 AVDD.t372 6.64567
R756 AVDD.n929 AVDD.t666 6.64567
R757 AVDD.n992 AVDD.t741 6.64567
R758 AVDD.n988 AVDD.t263 6.64567
R759 AVDD.n960 AVDD.t12 6.64567
R760 AVDD.n939 AVDD.t931 6.64567
R761 AVDD.n937 AVDD.t897 6.64567
R762 AVDD.n1048 AVDD.t1149 6.64567
R763 AVDD.n900 AVDD.t805 6.64567
R764 AVDD.n927 AVDD.t387 6.64567
R765 AVDD.n1753 AVDD.t1583 6.58663
R766 AVDD.n1703 AVDD.t1484 6.58663
R767 AVDD.n145 AVDD.t1358 6.58663
R768 AVDD.n232 AVDD.t1515 6.58663
R769 AVDD.n1916 AVDD.n1912 6.50088
R770 AVDD.n1865 AVDD.n1864 6.50088
R771 AVDD.n1587 AVDD.n1586 6.50088
R772 AVDD.n1540 AVDD.n1536 6.50088
R773 AVDD.n1708 AVDD.n1707 6.45575
R774 AVDD.n1659 AVDD.n1653 6.45575
R775 AVDD.n254 AVDD.n247 6.45575
R776 AVDD.n211 AVDD.n204 6.45575
R777 AVDD.n1754 AVDD.n1751 5.95439
R778 AVDD.n1704 AVDD.n1701 5.95439
R779 AVDD.n291 AVDD.n290 5.95439
R780 AVDD.n234 AVDD.n233 5.95439
R781 AVDD.n1751 AVDD.t1394 5.31528
R782 AVDD.n1701 AVDD.t1662 5.31528
R783 AVDD.n291 AVDD.t1555 5.31528
R784 AVDD.n234 AVDD.t1631 5.31528
R785 AVDD.n987 AVDD.t1379 5.19255
R786 AVDD.n1130 AVDD.t1414 5.12594
R787 AVDD.n1409 AVDD.n106 5.12014
R788 AVDD.n1951 AVDD.n37 5.12014
R789 AVDD.n951 AVDD.t1685 5.09041
R790 AVDD.t329 AVDD.n963 5.0505
R791 AVDD.n969 AVDD.t1184 5.0505
R792 AVDD.t992 AVDD.n970 5.0505
R793 AVDD.n971 AVDD.t992 5.0505
R794 AVDD.t265 AVDD.n989 5.0505
R795 AVDD.n995 AVDD.t667 5.0505
R796 AVDD.n1650 AVDD.n1649 4.96877
R797 AVDD.n1644 AVDD.n1643 4.96877
R798 AVDD.n208 AVDD.n207 4.96877
R799 AVDD.n251 AVDD.n250 4.96877
R800 AVDD.n49 AVDD.n47 4.92758
R801 AVDD.n1869 AVDD.n1867 4.92758
R802 AVDD.n72 AVDD.n70 4.92758
R803 AVDD.n1546 AVDD.n1544 4.92758
R804 AVDD.n1794 AVDD.n1793 4.78594
R805 AVDD.n1813 AVDD.n1812 4.78594
R806 AVDD.n1459 AVDD.n1458 4.78594
R807 AVDD.n1496 AVDD.n1495 4.78594
R808 AVDD.n1651 AVDD.n1650 4.61712
R809 AVDD.n1663 AVDD.n1662 4.61712
R810 AVDD.n1645 AVDD.n1644 4.61712
R811 AVDD.n1712 AVDD.n1711 4.61712
R812 AVDD.n209 AVDD.n208 4.61712
R813 AVDD.n199 AVDD.n198 4.61712
R814 AVDD.n252 AVDD.n251 4.61712
R815 AVDD.n242 AVDD.n241 4.61712
R816 AVDD.n1904 AVDD.n1901 4.61078
R817 AVDD.n1899 AVDD.n1896 4.61078
R818 AVDD.n1894 AVDD.n1891 4.61078
R819 AVDD.n1889 AVDD.n1886 4.61078
R820 AVDD.n1807 AVDD.n1804 4.61078
R821 AVDD.n1802 AVDD.n1799 4.61078
R822 AVDD.n1797 AVDD.n1794 4.61078
R823 AVDD.n1856 AVDD.n1853 4.61078
R824 AVDD.n1851 AVDD.n1848 4.61078
R825 AVDD.n1846 AVDD.n1843 4.61078
R826 AVDD.n1841 AVDD.n1838 4.61078
R827 AVDD.n1826 AVDD.n1823 4.61078
R828 AVDD.n1821 AVDD.n1818 4.61078
R829 AVDD.n1816 AVDD.n1813 4.61078
R830 AVDD.n1661 AVDD.n1660 4.61078
R831 AVDD.n1710 AVDD.n1709 4.61078
R832 AVDD.n1564 AVDD.n1563 4.61078
R833 AVDD.n1567 AVDD.n1566 4.61078
R834 AVDD.n1570 AVDD.n1569 4.61078
R835 AVDD.n1573 AVDD.n1572 4.61078
R836 AVDD.n1472 AVDD.n1469 4.61078
R837 AVDD.n1467 AVDD.n1464 4.61078
R838 AVDD.n1462 AVDD.n1459 4.61078
R839 AVDD.n1524 AVDD.n1523 4.61078
R840 AVDD.n1527 AVDD.n1526 4.61078
R841 AVDD.n1530 AVDD.n1529 4.61078
R842 AVDD.n1533 AVDD.n1532 4.61078
R843 AVDD.n1509 AVDD.n1506 4.61078
R844 AVDD.n1504 AVDD.n1501 4.61078
R845 AVDD.n1499 AVDD.n1496 4.61078
R846 AVDD.n203 AVDD.n200 4.61078
R847 AVDD.n246 AVDD.n243 4.61078
R848 AVDD.n1094 AVDD.n1090 4.61078
R849 AVDD.n1088 AVDD.n1084 4.61078
R850 AVDD.n1082 AVDD.n1078 4.61078
R851 AVDD.n1076 AVDD.n1074 4.61078
R852 AVDD.n1072 AVDD.n1068 4.61078
R853 AVDD.n1066 AVDD.n1062 4.61078
R854 AVDD.n1031 AVDD.n1030 4.61078
R855 AVDD.n1034 AVDD.n1033 4.61078
R856 AVDD.n1037 AVDD.n1036 4.61078
R857 AVDD.n1040 AVDD.n1039 4.61078
R858 AVDD.n1043 AVDD.n1042 4.61078
R859 AVDD.n1046 AVDD.n1045 4.61078
R860 AVDD.n1102 AVDD.n1101 4.60951
R861 AVDD.n1101 AVDD.n1100 4.60951
R862 AVDD.n1105 AVDD.n1104 4.60951
R863 AVDD.n1104 AVDD.n1103 4.60951
R864 AVDD.n1108 AVDD.n1107 4.60951
R865 AVDD.n1107 AVDD.n1106 4.60951
R866 AVDD.n1111 AVDD.n1110 4.60951
R867 AVDD.n1110 AVDD.n1109 4.60951
R868 AVDD.n1114 AVDD.n1113 4.60951
R869 AVDD.n1113 AVDD.n1112 4.60951
R870 AVDD.n1117 AVDD.n1116 4.60951
R871 AVDD.n1116 AVDD.n1115 4.60951
R872 AVDD.n1905 AVDD.n1904 4.60825
R873 AVDD.n1900 AVDD.n1899 4.60825
R874 AVDD.n1895 AVDD.n1894 4.60825
R875 AVDD.n1890 AVDD.n1889 4.60825
R876 AVDD.n1808 AVDD.n1807 4.60825
R877 AVDD.n1803 AVDD.n1802 4.60825
R878 AVDD.n1798 AVDD.n1797 4.60825
R879 AVDD.n1857 AVDD.n1856 4.60825
R880 AVDD.n1852 AVDD.n1851 4.60825
R881 AVDD.n1847 AVDD.n1846 4.60825
R882 AVDD.n1842 AVDD.n1841 4.60825
R883 AVDD.n1827 AVDD.n1826 4.60825
R884 AVDD.n1822 AVDD.n1821 4.60825
R885 AVDD.n1817 AVDD.n1816 4.60825
R886 AVDD.n1660 AVDD.n1659 4.60825
R887 AVDD.n1709 AVDD.n1708 4.60825
R888 AVDD.n1563 AVDD.n1562 4.60825
R889 AVDD.n1566 AVDD.n1565 4.60825
R890 AVDD.n1569 AVDD.n1568 4.60825
R891 AVDD.n1572 AVDD.n1571 4.60825
R892 AVDD.n1473 AVDD.n1472 4.60825
R893 AVDD.n1468 AVDD.n1467 4.60825
R894 AVDD.n1463 AVDD.n1462 4.60825
R895 AVDD.n1523 AVDD.n1486 4.60825
R896 AVDD.n1526 AVDD.n1525 4.60825
R897 AVDD.n1529 AVDD.n1528 4.60825
R898 AVDD.n1532 AVDD.n1531 4.60825
R899 AVDD.n1510 AVDD.n1509 4.60825
R900 AVDD.n1505 AVDD.n1504 4.60825
R901 AVDD.n1500 AVDD.n1499 4.60825
R902 AVDD.n204 AVDD.n203 4.60825
R903 AVDD.n247 AVDD.n246 4.60825
R904 AVDD.n1095 AVDD.n1094 4.60825
R905 AVDD.n1089 AVDD.n1088 4.60825
R906 AVDD.n1083 AVDD.n1082 4.60825
R907 AVDD.n1077 AVDD.n1076 4.60825
R908 AVDD.n1073 AVDD.n1072 4.60825
R909 AVDD.n1067 AVDD.n1066 4.60825
R910 AVDD.n1030 AVDD.n1029 4.60825
R911 AVDD.n1033 AVDD.n1032 4.60825
R912 AVDD.n1036 AVDD.n1035 4.60825
R913 AVDD.n1039 AVDD.n1038 4.60825
R914 AVDD.n1042 AVDD.n1041 4.60825
R915 AVDD.n1045 AVDD.n1044 4.60825
R916 AVDD.n1652 AVDD.n1651 4.60191
R917 AVDD.n1664 AVDD.n1663 4.60191
R918 AVDD.n1646 AVDD.n1645 4.60191
R919 AVDD.n1713 AVDD.n1712 4.60191
R920 AVDD.n210 AVDD.n209 4.60191
R921 AVDD.n198 AVDD.n179 4.60191
R922 AVDD.n253 AVDD.n252 4.60191
R923 AVDD.n241 AVDD.n239 4.60191
R924 AVDD.n1750 AVDD.n1748 4.50663
R925 AVDD.n1700 AVDD.n1635 4.50663
R926 AVDD.n294 AVDD.n293 4.50663
R927 AVDD.n237 AVDD.n236 4.50663
R928 AVDD.n1796 AVDD.n1792 4.5005
R929 AVDD.n1801 AVDD.n1791 4.5005
R930 AVDD.n1806 AVDD.n1790 4.5005
R931 AVDD.n1888 AVDD.n1789 4.5005
R932 AVDD.n1893 AVDD.n1788 4.5005
R933 AVDD.n1898 AVDD.n1787 4.5005
R934 AVDD.n1903 AVDD.n1786 4.5005
R935 AVDD.n1815 AVDD.n1811 4.5005
R936 AVDD.n1820 AVDD.n1810 4.5005
R937 AVDD.n1825 AVDD.n1809 4.5005
R938 AVDD.n1840 AVDD.n1837 4.5005
R939 AVDD.n1845 AVDD.n1836 4.5005
R940 AVDD.n1850 AVDD.n1835 4.5005
R941 AVDD.n1855 AVDD.n1834 4.5005
R942 AVDD.n1637 AVDD.n1636 4.5005
R943 AVDD.n1640 AVDD.n1638 4.5005
R944 AVDD.n1642 AVDD.n1641 4.5005
R945 AVDD.n1655 AVDD.n1654 4.5005
R946 AVDD.n1658 AVDD.n1656 4.5005
R947 AVDD.n1648 AVDD.n1647 4.5005
R948 AVDD.n1461 AVDD.n1457 4.5005
R949 AVDD.n1466 AVDD.n1456 4.5005
R950 AVDD.n1471 AVDD.n1455 4.5005
R951 AVDD.n1476 AVDD.n1474 4.5005
R952 AVDD.n1479 AVDD.n1477 4.5005
R953 AVDD.n1482 AVDD.n1480 4.5005
R954 AVDD.n1485 AVDD.n1483 4.5005
R955 AVDD.n1498 AVDD.n1494 4.5005
R956 AVDD.n1503 AVDD.n1493 4.5005
R957 AVDD.n1508 AVDD.n1492 4.5005
R958 AVDD.n1513 AVDD.n1511 4.5005
R959 AVDD.n1516 AVDD.n1514 4.5005
R960 AVDD.n1519 AVDD.n1517 4.5005
R961 AVDD.n1522 AVDD.n1520 4.5005
R962 AVDD.n240 AVDD.n178 4.5005
R963 AVDD.n245 AVDD.n177 4.5005
R964 AVDD.n249 AVDD.n248 4.5005
R965 AVDD.n197 AVDD.n196 4.5005
R966 AVDD.n202 AVDD.n195 4.5005
R967 AVDD.n206 AVDD.n205 4.5005
R968 AVDD.n668 AVDD.n666 4.5005
R969 AVDD.n671 AVDD.n669 4.5005
R970 AVDD.n673 AVDD.n672 4.5005
R971 AVDD.n676 AVDD.n674 4.5005
R972 AVDD.n679 AVDD.n677 4.5005
R973 AVDD.n682 AVDD.n680 4.5005
R974 AVDD.n1064 AVDD.n692 4.5005
R975 AVDD.n1070 AVDD.n691 4.5005
R976 AVDD.n1075 AVDD.n690 4.5005
R977 AVDD.n1080 AVDD.n689 4.5005
R978 AVDD.n1086 AVDD.n688 4.5005
R979 AVDD.n1092 AVDD.n687 4.5005
R980 AVDD.n903 AVDD.n901 4.5005
R981 AVDD.n906 AVDD.n904 4.5005
R982 AVDD.n908 AVDD.n907 4.5005
R983 AVDD.n911 AVDD.n909 4.5005
R984 AVDD.n914 AVDD.n912 4.5005
R985 AVDD.n917 AVDD.n915 4.5005
R986 AVDD.n1665 AVDD.n1664 4.32507
R987 AVDD.n230 AVDD.n179 4.32507
R988 AVDD.n1859 AVDD.t1392 4.06712
R989 AVDD.n1832 AVDD.t1292 4.06712
R990 AVDD.n1917 AVDD.t1683 4.06712
R991 AVDD.n1910 AVDD.t1408 4.06712
R992 AVDD.n1541 AVDD.t1377 4.06712
R993 AVDD.n1490 AVDD.t1504 4.06712
R994 AVDD.n1581 AVDD.t1373 4.06712
R995 AVDD.n1579 AVDD.t1348 4.06712
R996 AVDD.n1919 AVDD.n1918 3.96014
R997 AVDD.n1860 AVDD.n1858 3.96014
R998 AVDD.n1582 AVDD.n69 3.96014
R999 AVDD.n1543 AVDD.n1542 3.96014
R1000 AVDD.n1859 AVDD.t1422 3.86107
R1001 AVDD.n1832 AVDD.t1453 3.86107
R1002 AVDD.n1917 AVDD.t1594 3.86107
R1003 AVDD.n1910 AVDD.t1401 3.86107
R1004 AVDD.n1541 AVDD.t1346 3.86107
R1005 AVDD.n1490 AVDD.t1623 3.86107
R1006 AVDD.n1581 AVDD.t1363 3.86107
R1007 AVDD.n1579 AVDD.t1562 3.86107
R1008 AVDD.n1648 AVDD.t1588 3.84568
R1009 AVDD.n1655 AVDD.t1300 3.84568
R1010 AVDD.n1642 AVDD.t1567 3.84568
R1011 AVDD.n1637 AVDD.t1686 3.84568
R1012 AVDD.n206 AVDD.t1333 3.84568
R1013 AVDD.n197 AVDD.t1537 3.84568
R1014 AVDD.n249 AVDD.t1611 3.84568
R1015 AVDD.n240 AVDD.t1318 3.84568
R1016 AVDD.n1753 AVDD.n1752 3.84528
R1017 AVDD.n1750 AVDD.n1749 3.84528
R1018 AVDD.n1703 AVDD.n1702 3.84528
R1019 AVDD.n1700 AVDD.n1699 3.84528
R1020 AVDD.n145 AVDD.n144 3.84528
R1021 AVDD.n293 AVDD.n292 3.84528
R1022 AVDD.n232 AVDD.n231 3.84528
R1023 AVDD.n236 AVDD.n235 3.84528
R1024 AVDD.n1076 AVDD.t1694 3.84449
R1025 AVDD.n51 AVDD.n49 3.79678
R1026 AVDD.n1926 AVDD.n1924 3.79678
R1027 AVDD.n1871 AVDD.n1869 3.79678
R1028 AVDD.n1879 AVDD.n1877 3.79678
R1029 AVDD.n1742 AVDD.n1738 3.79678
R1030 AVDD.n1725 AVDD.n1721 3.79678
R1031 AVDD.n1677 AVDD.n1673 3.79678
R1032 AVDD.n1692 AVDD.n1688 3.79678
R1033 AVDD.n74 AVDD.n72 3.79678
R1034 AVDD.n1596 AVDD.n1594 3.79678
R1035 AVDD.n1548 AVDD.n1546 3.79678
R1036 AVDD.n1557 AVDD.n1555 3.79678
R1037 AVDD.n267 AVDD.n263 3.79678
R1038 AVDD.n282 AVDD.n278 3.79678
R1039 AVDD.n225 AVDD.n221 3.79678
R1040 AVDD.n190 AVDD.n186 3.79678
R1041 AVDD.n1714 AVDD.n1713 3.74038
R1042 AVDD.n239 AVDD.n238 3.74038
R1043 AVDD.n1734 AVDD.n1730 3.73034
R1044 AVDD.n1697 AVDD.n1681 3.73034
R1045 AVDD.n287 AVDD.n271 3.73034
R1046 AVDD.n217 AVDD.n213 3.73034
R1047 AVDD.n1055 AVDD.t717 3.7109
R1048 AVDD.n1075 AVDD.t1282 3.68344
R1049 AVDD.n1129 AVDD.n1128 3.65594
R1050 AVDD.n1922 AVDD.n1921 3.65581
R1051 AVDD.n1924 AVDD.n1923 3.65581
R1052 AVDD.n1926 AVDD.n1925 3.65581
R1053 AVDD.n1928 AVDD.n1927 3.65581
R1054 AVDD.n53 AVDD.n52 3.65581
R1055 AVDD.n51 AVDD.n50 3.65581
R1056 AVDD.n49 AVDD.n48 3.65581
R1057 AVDD.n1875 AVDD.n1874 3.65581
R1058 AVDD.n1877 AVDD.n1876 3.65581
R1059 AVDD.n1879 AVDD.n1878 3.65581
R1060 AVDD.n1881 AVDD.n1880 3.65581
R1061 AVDD.n1873 AVDD.n1872 3.65581
R1062 AVDD.n1871 AVDD.n1870 3.65581
R1063 AVDD.n1869 AVDD.n1868 3.65581
R1064 AVDD.n1598 AVDD.n1597 3.65581
R1065 AVDD.n1596 AVDD.n1595 3.65581
R1066 AVDD.n1594 AVDD.n1593 3.65581
R1067 AVDD.n1592 AVDD.n1591 3.65581
R1068 AVDD.n76 AVDD.n75 3.65581
R1069 AVDD.n74 AVDD.n73 3.65581
R1070 AVDD.n72 AVDD.n71 3.65581
R1071 AVDD.n1559 AVDD.n1558 3.65581
R1072 AVDD.n1557 AVDD.n1556 3.65581
R1073 AVDD.n1555 AVDD.n1554 3.65581
R1074 AVDD.n1553 AVDD.n1552 3.65581
R1075 AVDD.n1550 AVDD.n1549 3.65581
R1076 AVDD.n1548 AVDD.n1547 3.65581
R1077 AVDD.n1546 AVDD.n1545 3.65581
R1078 AVDD.n1134 AVDD.n1133 3.6512
R1079 AVDD.n1125 AVDD.n1124 3.6512
R1080 AVDD.n1132 AVDD.n1131 3.6512
R1081 AVDD.n1127 AVDD.n1126 3.6512
R1082 AVDD.n1929 AVDD.n1928 3.64443
R1083 AVDD.n1882 AVDD.n1881 3.64443
R1084 AVDD.n1592 AVDD.n1590 3.64443
R1085 AVDD.n1553 AVDD.n1551 3.64443
R1086 AVDD.n908 AVDD.t1427 3.6266
R1087 AVDD.n948 AVDD.n947 3.62041
R1088 AVDD.n950 AVDD.n949 3.62041
R1089 AVDD.n953 AVDD.n952 3.62041
R1090 AVDD.n955 AVDD.n954 3.62041
R1091 AVDD.n957 AVDD.n956 3.62041
R1092 AVDD.n673 AVDD.t1663 3.61594
R1093 AVDD.n1799 AVDD.n1798 3.524
R1094 AVDD.n1896 AVDD.n1895 3.524
R1095 AVDD.n1818 AVDD.n1817 3.524
R1096 AVDD.n1848 AVDD.n1847 3.524
R1097 AVDD.n1464 AVDD.n1463 3.524
R1098 AVDD.n1568 AVDD.n1567 3.524
R1099 AVDD.n1501 AVDD.n1500 3.524
R1100 AVDD.n1528 AVDD.n1527 3.524
R1101 AVDD.n1886 AVDD.n1885 3.506
R1102 AVDD.n1838 AVDD.n1828 3.506
R1103 AVDD.n1574 AVDD.n1573 3.506
R1104 AVDD.n1534 AVDD.n1533 3.506
R1105 AVDD.n1604 AVDD.t139 3.20383
R1106 AVDD.n158 AVDD.t422 3.20383
R1107 AVDD.t384 AVDD.n159 3.20383
R1108 AVDD.n166 AVDD.t1076 3.20383
R1109 AVDD.t1108 AVDD.n167 3.20383
R1110 AVDD.t934 AVDD.n148 3.20383
R1111 AVDD.n1935 AVDD.t1208 3.20383
R1112 AVDD.n1617 AVDD.t1064 3.20383
R1113 AVDD.t1136 AVDD.n1618 3.20383
R1114 AVDD.n1625 AVDD.t418 3.20383
R1115 AVDD.t287 AVDD.n1626 3.20383
R1116 AVDD.t1168 AVDD.n1607 3.20383
R1117 AVDD.t105 AVDD.n1227 3.20383
R1118 AVDD.n1228 AVDD.t105 3.20383
R1119 AVDD.n1229 AVDD.t665 3.20383
R1120 AVDD.n1238 AVDD.t904 3.20383
R1121 AVDD.t527 AVDD.n1239 3.20383
R1122 AVDD.n1246 AVDD.t501 3.20383
R1123 AVDD.n1247 AVDD.t91 3.20383
R1124 AVDD.n1256 AVDD.t1098 3.20383
R1125 AVDD.t9 AVDD.n1257 3.20383
R1126 AVDD.n1258 AVDD.t9 3.20383
R1127 AVDD.t938 AVDD.n1263 3.20383
R1128 AVDD.n1264 AVDD.t938 3.20383
R1129 AVDD.n1265 AVDD.t1158 3.20383
R1130 AVDD.n1274 AVDD.t426 3.20383
R1131 AVDD.t1016 AVDD.n1275 3.20383
R1132 AVDD.n1282 AVDD.t6 3.20383
R1133 AVDD.n1283 AVDD.t594 3.20383
R1134 AVDD.n1292 AVDD.t1210 3.20383
R1135 AVDD.n1227 AVDD.t117 3.20383
R1136 AVDD.n1228 AVDD.t117 3.20383
R1137 AVDD.n1229 AVDD.t673 3.20383
R1138 AVDD.n1238 AVDD.t910 3.20383
R1139 AVDD.n1239 AVDD.t533 3.20383
R1140 AVDD.n1246 AVDD.t509 3.20383
R1141 AVDD.n1247 AVDD.t103 3.20383
R1142 AVDD.n1256 AVDD.t1104 3.20383
R1143 AVDD.n1257 AVDD.t25 3.20383
R1144 AVDD.n1258 AVDD.t25 3.20383
R1145 AVDD.n1263 AVDD.t942 3.20383
R1146 AVDD.n1264 AVDD.t942 3.20383
R1147 AVDD.n1265 AVDD.t1166 3.20383
R1148 AVDD.n1274 AVDD.t430 3.20383
R1149 AVDD.n1275 AVDD.t1020 3.20383
R1150 AVDD.n1282 AVDD.t11 3.20383
R1151 AVDD.n1283 AVDD.t600 3.20383
R1152 AVDD.n1292 AVDD.t1216 3.20383
R1153 AVDD.n1203 AVDD.t1246 3.20383
R1154 AVDD.t1246 AVDD.n1202 3.20383
R1155 AVDD.n1201 AVDD.t715 3.20383
R1156 AVDD.n1191 AVDD.t900 3.20383
R1157 AVDD.n1190 AVDD.t620 3.20383
R1158 AVDD.t239 AVDD.n1183 3.20383
R1159 AVDD.n1182 AVDD.t489 3.20383
R1160 AVDD.t206 AVDD.n32 3.20383
R1161 AVDD.n1782 AVDD.t819 3.20383
R1162 AVDD.n1773 AVDD.t996 3.20383
R1163 AVDD.n1772 AVDD.t732 3.20383
R1164 AVDD.t343 AVDD.n1765 3.20383
R1165 AVDD.n1764 AVDD.t586 3.20383
R1166 AVDD.t311 AVDD.n42 3.20383
R1167 AVDD.n1961 AVDD.t1112 3.20383
R1168 AVDD.n1970 AVDD.t988 3.20383
R1169 AVDD.t1024 AVDD.n1971 3.20383
R1170 AVDD.n1301 AVDD.t331 3.20383
R1171 AVDD.n1302 AVDD.t154 3.20383
R1172 AVDD.n1311 AVDD.t1056 3.20383
R1173 AVDD.n1961 AVDD.t466 3.20383
R1174 AVDD.n1970 AVDD.t341 3.20383
R1175 AVDD.n1971 AVDD.t376 3.20383
R1176 AVDD.n1301 AVDD.t964 3.20383
R1177 AVDD.n1302 AVDD.t813 3.20383
R1178 AVDD.n1311 AVDD.t412 3.20383
R1179 AVDD.n501 AVDD.t736 3.20383
R1180 AVDD.n491 AVDD.t699 3.20383
R1181 AVDD.n490 AVDD.t970 3.20383
R1182 AVDD.t382 AVDD.n483 3.20383
R1183 AVDD.n482 AVDD.t348 3.20383
R1184 AVDD.n472 AVDD.t1200 3.20383
R1185 AVDD.n471 AVDD.t151 3.20383
R1186 AVDD.t151 AVDD.n470 3.20383
R1187 AVDD.n501 AVDD.t1140 3.20383
R1188 AVDD.t1078 AVDD.n491 3.20383
R1189 AVDD.n490 AVDD.t60 3.20383
R1190 AVDD.n483 AVDD.t804 3.20383
R1191 AVDD.n482 AVDD.t758 3.20383
R1192 AVDD.t333 AVDD.n472 3.20383
R1193 AVDD.n471 AVDD.t570 3.20383
R1194 AVDD.n470 AVDD.t570 3.20383
R1195 AVDD.t558 AVDD.n12 3.20383
R1196 AVDD.n419 AVDD.t839 3.20383
R1197 AVDD.t796 AVDD.n420 3.20383
R1198 AVDD.n427 AVDD.t201 3.20383
R1199 AVDD.n428 AVDD.t227 3.20383
R1200 AVDD.n437 AVDD.t1280 3.20383
R1201 AVDD.t950 AVDD.n12 3.20383
R1202 AVDD.n419 AVDD.t1218 3.20383
R1203 AVDD.n420 AVDD.t1176 3.20383
R1204 AVDD.n427 AVDD.t612 3.20383
R1205 AVDD.n428 AVDD.t630 3.20383
R1206 AVDD.n437 AVDD.t434 3.20383
R1207 AVDD.n1378 AVDD.t454 3.20383
R1208 AVDD.n1387 AVDD.t762 3.20383
R1209 AVDD.t157 AVDD.n1388 3.20383
R1210 AVDD.t1146 AVDD.n613 3.20383
R1211 AVDD.n610 AVDD.t462 3.20383
R1212 AVDD.n600 AVDD.t244 3.20383
R1213 AVDD.n599 AVDD.t968 3.20383
R1214 AVDD.t968 AVDD.n598 3.20383
R1215 AVDD.n596 AVDD.t408 3.20383
R1216 AVDD.t408 AVDD.n595 3.20383
R1217 AVDD.n594 AVDD.t1148 3.20383
R1218 AVDD.n584 AVDD.t460 3.20383
R1219 AVDD.n583 AVDD.t859 3.20383
R1220 AVDD.t531 AVDD.n576 3.20383
R1221 AVDD.n575 AVDD.t1224 3.20383
R1222 AVDD.n565 AVDD.t821 3.20383
R1223 AVDD.n564 AVDD.t592 3.20383
R1224 AVDD.t592 AVDD.n563 3.20383
R1225 AVDD.n1378 AVDD.t464 3.20383
R1226 AVDD.n1387 AVDD.t770 3.20383
R1227 AVDD.n1388 AVDD.t161 3.20383
R1228 AVDD.n613 AVDD.t1152 3.20383
R1229 AVDD.n610 AVDD.t474 3.20383
R1230 AVDD.t250 AVDD.n600 3.20383
R1231 AVDD.n599 AVDD.t976 3.20383
R1232 AVDD.n598 AVDD.t976 3.20383
R1233 AVDD.n596 AVDD.t410 3.20383
R1234 AVDD.n595 AVDD.t410 3.20383
R1235 AVDD.n594 AVDD.t1156 3.20383
R1236 AVDD.t468 AVDD.n584 3.20383
R1237 AVDD.n583 AVDD.t861 3.20383
R1238 AVDD.n576 AVDD.t539 3.20383
R1239 AVDD.n575 AVDD.t1230 3.20383
R1240 AVDD.t829 AVDD.n565 3.20383
R1241 AVDD.n564 AVDD.t598 3.20383
R1242 AVDD.n563 AVDD.t598 3.20383
R1243 AVDD.n518 AVDD.t275 3.20383
R1244 AVDD.n527 AVDD.t218 3.20383
R1245 AVDD.t491 AVDD.n528 3.20383
R1246 AVDD.n535 AVDD.t1190 3.20383
R1247 AVDD.n536 AVDD.t1160 3.20383
R1248 AVDD.n545 AVDD.t750 3.20383
R1249 AVDD.t51 AVDD.n15 3.20383
R1250 AVDD.n378 AVDD.t360 3.20383
R1251 AVDD.t317 AVDD.n379 3.20383
R1252 AVDD.n386 AVDD.t1012 3.20383
R1253 AVDD.n387 AVDD.t1028 3.20383
R1254 AVDD.n396 AVDD.t873 3.20383
R1255 AVDD.n1419 AVDD.t242 3.20383
R1256 AVDD.n1428 AVDD.t194 3.20383
R1257 AVDD.t456 AVDD.n1429 3.20383
R1258 AVDD.n331 AVDD.t1172 3.20383
R1259 AVDD.n332 AVDD.t1128 3.20383
R1260 AVDD.n341 AVDD.t728 3.20383
R1261 AVDD.n342 AVDD.t952 3.20383
R1262 AVDD.t952 AVDD.n322 3.20383
R1263 AVDD.n1419 AVDD.t886 3.20383
R1264 AVDD.n1428 AVDD.t847 3.20383
R1265 AVDD.n1429 AVDD.t1092 3.20383
R1266 AVDD.n331 AVDD.t525 3.20383
R1267 AVDD.n332 AVDD.t483 3.20383
R1268 AVDD.n341 AVDD.t45 3.20383
R1269 AVDD.n342 AVDD.t309 3.20383
R1270 AVDD.t309 AVDD.n322 3.20383
R1271 AVDD.n1451 AVDD.t345 3.20383
R1272 AVDD.n1442 AVDD.t307 3.20383
R1273 AVDD.n1441 AVDD.t576 3.20383
R1274 AVDD.n299 AVDD.t1254 3.20383
R1275 AVDD.n300 AVDD.t1214 3.20383
R1276 AVDD.n309 AVDD.t827 3.20383
R1277 AVDD.n1351 AVDD.t23 3.20383
R1278 AVDD.n1341 AVDD.t339 3.20383
R1279 AVDD.n1340 AVDD.t299 3.20383
R1280 AVDD.t994 AVDD.n1333 3.20383
R1281 AVDD.n1332 AVDD.t1010 3.20383
R1282 AVDD.t845 AVDD.n101 3.20383
R1283 AVDD.n1351 AVDD.t693 3.20383
R1284 AVDD.t974 AVDD.n1341 3.20383
R1285 AVDD.n1340 AVDD.t928 3.20383
R1286 AVDD.n1333 AVDD.t352 3.20383
R1287 AVDD.n1332 AVDD.t369 3.20383
R1288 AVDD.t179 AVDD.n101 3.20383
R1289 AVDD.n710 AVDD.t922 3.20383
R1290 AVDD.n707 AVDD.t641 3.20383
R1291 AVDD.t273 AVDD.n703 3.20383
R1292 AVDD.n699 AVDD.t511 3.20383
R1293 AVDD.t229 AVDD.n881 3.20383
R1294 AVDD.n877 AVDD.t1250 3.20383
R1295 AVDD.t1250 AVDD.n876 3.20383
R1296 AVDD.n870 AVDD.t77 3.20383
R1297 AVDD.t77 AVDD.n869 3.20383
R1298 AVDD.n866 AVDD.t1154 3.20383
R1299 AVDD.t655 AVDD.n661 3.20383
R1300 AVDD.n662 AVDD.t655 3.20383
R1301 AVDD.t1204 AVDD.n712 3.20383
R1302 AVDD.n723 AVDD.t1252 3.20383
R1303 AVDD.n887 AVDD.t1044 3.20383
R1304 AVDD.t28 AVDD.n884 3.20383
R1305 AVDD.n880 AVDD.t687 3.20383
R1306 AVDD.n867 AVDD.t476 3.20383
R1307 AVDD.t616 AVDD.n848 3.20383
R1308 AVDD.n858 AVDD.t616 3.20383
R1309 AVDD.n1146 AVDD.t740 3.20383
R1310 AVDD.t1006 AVDD.n854 3.20383
R1311 AVDD.n853 AVDD.t1042 3.20383
R1312 AVDD.n1982 AVDD.t356 3.20383
R1313 AVDD.n1983 AVDD.t184 3.20383
R1314 AVDD.n1992 AVDD.t1074 3.20383
R1315 AVDD.n821 AVDD.t336 3.20383
R1316 AVDD.n811 AVDD.t196 3.20383
R1317 AVDD.n810 AVDD.t253 3.20383
R1318 AVDD.t835 AVDD.n803 3.20383
R1319 AVDD.n802 AVDD.t663 3.20383
R1320 AVDD.t295 AVDD.n13 3.20383
R1321 AVDD.n821 AVDD.t746 3.20383
R1322 AVDD.t602 AVDD.n811 3.20383
R1323 AVDD.n810 AVDD.t647 3.20383
R1324 AVDD.n803 AVDD.t1212 3.20383
R1325 AVDD.n802 AVDD.t1054 3.20383
R1326 AVDD.t683 AVDD.n13 3.20383
R1327 AVDD.t478 AVDD.n751 3.20383
R1328 AVDD.n752 AVDD.t478 3.20383
R1329 AVDD.n753 AVDD.t1198 3.20383
R1330 AVDD.n762 AVDD.t94 3.20383
R1331 AVDD.t1102 AVDD.n763 3.20383
R1332 AVDD.n770 AVDD.t734 3.20383
R1333 AVDD.n771 AVDD.t986 3.20383
R1334 AVDD.n780 AVDD.t709 3.20383
R1335 AVDD.n751 AVDD.t896 3.20383
R1336 AVDD.n752 AVDD.t896 3.20383
R1337 AVDD.n753 AVDD.t326 3.20383
R1338 AVDD.n762 AVDD.t507 3.20383
R1339 AVDD.n763 AVDD.t234 3.20383
R1340 AVDD.n770 AVDD.t1138 3.20383
R1341 AVDD.n771 AVDD.t83 3.20383
R1342 AVDD.n780 AVDD.t1088 3.20383
R1343 AVDD.n1025 AVDD.t811 3.20383
R1344 AVDD.n1016 AVDD.t876 3.20383
R1345 AVDD.n1015 AVDD.t639 3.20383
R1346 AVDD.t926 AVDD.n1008 3.20383
R1347 AVDD.n1007 AVDD.t283 3.20383
R1348 AVDD.n998 AVDD.t40 3.20383
R1349 AVDD.n1203 AVDD.t622 3.20383
R1350 AVDD.n1202 AVDD.t622 3.20383
R1351 AVDD.n1201 AVDD.t34 3.20383
R1352 AVDD.t258 AVDD.n1191 3.20383
R1353 AVDD.n1190 AVDD.t1240 3.20383
R1354 AVDD.n1183 AVDD.t884 3.20383
R1355 AVDD.n1182 AVDD.t1114 3.20383
R1356 AVDD.t851 AVDD.n32 3.20383
R1357 AVDD.n1754 AVDD.n1753 3.00663
R1358 AVDD.n1704 AVDD.n1703 3.00663
R1359 AVDD.n290 AVDD.n145 3.00663
R1360 AVDD.n233 AVDD.n232 3.00663
R1361 AVDD.n1717 AVDD.n1715 2.7866
R1362 AVDD.n1720 AVDD.n1718 2.7866
R1363 AVDD.n1724 AVDD.n1722 2.7866
R1364 AVDD.n1728 AVDD.n1726 2.7866
R1365 AVDD.n1733 AVDD.n1731 2.7866
R1366 AVDD.n1737 AVDD.n1735 2.7866
R1367 AVDD.n1741 AVDD.n1739 2.7866
R1368 AVDD.n1745 AVDD.n1743 2.7866
R1369 AVDD.n1684 AVDD.n1682 2.7866
R1370 AVDD.n1687 AVDD.n1685 2.7866
R1371 AVDD.n1691 AVDD.n1689 2.7866
R1372 AVDD.n1695 AVDD.n1693 2.7866
R1373 AVDD.n1680 AVDD.n1678 2.7866
R1374 AVDD.n1676 AVDD.n1674 2.7866
R1375 AVDD.n1672 AVDD.n1670 2.7866
R1376 AVDD.n1668 AVDD.n1666 2.7866
R1377 AVDD.n274 AVDD.n272 2.7866
R1378 AVDD.n277 AVDD.n275 2.7866
R1379 AVDD.n281 AVDD.n279 2.7866
R1380 AVDD.n285 AVDD.n283 2.7866
R1381 AVDD.n270 AVDD.n268 2.7866
R1382 AVDD.n266 AVDD.n264 2.7866
R1383 AVDD.n262 AVDD.n260 2.7866
R1384 AVDD.n258 AVDD.n256 2.7866
R1385 AVDD.n182 AVDD.n180 2.7866
R1386 AVDD.n185 AVDD.n183 2.7866
R1387 AVDD.n189 AVDD.n187 2.7866
R1388 AVDD.n193 AVDD.n191 2.7866
R1389 AVDD.n216 AVDD.n214 2.7866
R1390 AVDD.n220 AVDD.n218 2.7866
R1391 AVDD.n224 AVDD.n222 2.7866
R1392 AVDD.n228 AVDD.n226 2.7866
R1393 AVDD.n1911 AVDD.n1909 2.73714
R1394 AVDD.n1833 AVDD.n1831 2.73714
R1395 AVDD.n1580 AVDD.n1578 2.73714
R1396 AVDD.n1491 AVDD.n1489 2.73714
R1397 AVDD.n1721 AVDD.n1717 2.73672
R1398 AVDD.n1688 AVDD.n1684 2.73672
R1399 AVDD.n278 AVDD.n274 2.73672
R1400 AVDD.n186 AVDD.n182 2.73672
R1401 AVDD.n958 AVDD.n957 2.60496
R1402 AVDD.n1125 AVDD.n1123 2.60386
R1403 AVDD.n991 AVDD.n990 2.6005
R1404 AVDD.n994 AVDD.n993 2.6005
R1405 AVDD.n968 AVDD.n967 2.6005
R1406 AVDD.n965 AVDD.n964 2.6005
R1407 AVDD.n948 AVDD.n946 2.59852
R1408 AVDD.n1135 AVDD.n1134 2.59742
R1409 AVDD.n1863 AVDD.n1861 2.59712
R1410 AVDD.n1831 AVDD.n1829 2.59712
R1411 AVDD.n1915 AVDD.n1913 2.59712
R1412 AVDD.n1909 AVDD.n1907 2.59712
R1413 AVDD.n1539 AVDD.n1537 2.59712
R1414 AVDD.n1489 AVDD.n1487 2.59712
R1415 AVDD.n1585 AVDD.n1583 2.59712
R1416 AVDD.n1578 AVDD.n1576 2.59712
R1417 AVDD.n972 AVDD.t1276 2.5255
R1418 AVDD.n974 AVDD.t920 2.5255
R1419 AVDD.n977 AVDD.t543 2.5255
R1420 AVDD.n977 AVDD.t888 2.5255
R1421 AVDD.n981 AVDD.t808 2.5255
R1422 AVDD.n981 AVDD.t1132 2.5255
R1423 AVDD.n984 AVDD.t436 2.5255
R1424 AVDD.n984 AVDD.t798 2.5255
R1425 AVDD.n986 AVDD.t3 2.5255
R1426 AVDD.n986 AVDD.t374 2.5255
R1427 AVDD.n961 AVDD.t14 2.5255
R1428 AVDD.n940 AVDD.t932 2.5255
R1429 AVDD.n935 AVDD.t898 2.5255
R1430 AVDD.n1049 AVDD.t1150 2.5255
R1431 AVDD.n925 AVDD.t806 2.5255
R1432 AVDD.n996 AVDD.t388 2.5255
R1433 AVDD.n1118 AVDD.n1117 2.46986
R1434 AVDD.n1062 AVDD.n1061 2.46873
R1435 AVDD.n1047 AVDD.n1046 2.46873
R1436 AVDD.n1029 AVDD.n1028 2.46198
R1437 AVDD.n1096 AVDD.n1095 2.46198
R1438 AVDD.n1100 AVDD.n1099 2.46086
R1439 AVDD.n1912 AVDD.n1911 2.46014
R1440 AVDD.n1865 AVDD.n1833 2.46014
R1441 AVDD.n1587 AVDD.n1580 2.46014
R1442 AVDD.n1536 AVDD.n1491 2.46014
R1443 AVDD.n964 AVDD.t395 2.4505
R1444 AVDD.n964 AVDD.t329 2.4505
R1445 AVDD.t1184 AVDD.n968 2.4505
R1446 AVDD.n968 AVDD.t395 2.4505
R1447 AVDD.n994 AVDD.t742 2.4505
R1448 AVDD.t667 AVDD.n994 2.4505
R1449 AVDD.n990 AVDD.t265 2.4505
R1450 AVDD.n990 AVDD.t742 2.4505
R1451 AVDD.n1863 AVDD.n1862 2.39107
R1452 AVDD.n1831 AVDD.n1830 2.39107
R1453 AVDD.n1915 AVDD.n1914 2.39107
R1454 AVDD.n1909 AVDD.n1908 2.39107
R1455 AVDD.n1539 AVDD.n1538 2.39107
R1456 AVDD.n1489 AVDD.n1488 2.39107
R1457 AVDD.n1585 AVDD.n1584 2.39107
R1458 AVDD.n1578 AVDD.n1577 2.39107
R1459 AVDD.n1658 AVDD.n1657 2.37568
R1460 AVDD.n1640 AVDD.n1639 2.37568
R1461 AVDD.n202 AVDD.n201 2.37568
R1462 AVDD.n245 AVDD.n244 2.37568
R1463 AVDD.n1094 AVDD.n1093 2.37449
R1464 AVDD.n1088 AVDD.n1087 2.37449
R1465 AVDD.n1082 AVDD.n1081 2.37449
R1466 AVDD.n1072 AVDD.n1071 2.37449
R1467 AVDD.n1066 AVDD.n1065 2.37449
R1468 AVDD.n1931 AVDD.n43 2.30165
R1469 AVDD.n1784 AVDD.n1783 2.30165
R1470 AVDD.n1600 AVDD.n66 2.30165
R1471 AVDD.n1453 AVDD.n1452 2.30165
R1472 AVDD.n1707 AVDD.n1646 2.24038
R1473 AVDD.n1653 AVDD.n1652 2.24038
R1474 AVDD.n254 AVDD.n253 2.24038
R1475 AVDD.n211 AVDD.n210 2.24038
R1476 AVDD.n1092 AVDD.n1091 2.21344
R1477 AVDD.n1086 AVDD.n1085 2.21344
R1478 AVDD.n1080 AVDD.n1079 2.21344
R1479 AVDD.n1070 AVDD.n1069 2.21344
R1480 AVDD.n1064 AVDD.n1063 2.21344
R1481 AVDD.n1717 AVDD.n1716 2.2016
R1482 AVDD.n1720 AVDD.n1719 2.2016
R1483 AVDD.n1724 AVDD.n1723 2.2016
R1484 AVDD.n1728 AVDD.n1727 2.2016
R1485 AVDD.n1733 AVDD.n1732 2.2016
R1486 AVDD.n1737 AVDD.n1736 2.2016
R1487 AVDD.n1741 AVDD.n1740 2.2016
R1488 AVDD.n1745 AVDD.n1744 2.2016
R1489 AVDD.n1684 AVDD.n1683 2.2016
R1490 AVDD.n1687 AVDD.n1686 2.2016
R1491 AVDD.n1691 AVDD.n1690 2.2016
R1492 AVDD.n1695 AVDD.n1694 2.2016
R1493 AVDD.n1680 AVDD.n1679 2.2016
R1494 AVDD.n1676 AVDD.n1675 2.2016
R1495 AVDD.n1672 AVDD.n1671 2.2016
R1496 AVDD.n1668 AVDD.n1667 2.2016
R1497 AVDD.n274 AVDD.n273 2.2016
R1498 AVDD.n277 AVDD.n276 2.2016
R1499 AVDD.n281 AVDD.n280 2.2016
R1500 AVDD.n285 AVDD.n284 2.2016
R1501 AVDD.n270 AVDD.n269 2.2016
R1502 AVDD.n266 AVDD.n265 2.2016
R1503 AVDD.n262 AVDD.n261 2.2016
R1504 AVDD.n258 AVDD.n257 2.2016
R1505 AVDD.n182 AVDD.n181 2.2016
R1506 AVDD.n185 AVDD.n184 2.2016
R1507 AVDD.n189 AVDD.n188 2.2016
R1508 AVDD.n193 AVDD.n192 2.2016
R1509 AVDD.n216 AVDD.n215 2.2016
R1510 AVDD.n220 AVDD.n219 2.2016
R1511 AVDD.n224 AVDD.n223 2.2016
R1512 AVDD.n228 AVDD.n227 2.2016
R1513 AVDD.n1858 AVDD.n1857 2.18645
R1514 AVDD.n1543 AVDD.n1486 2.18645
R1515 AVDD.n1903 AVDD.n1902 2.18502
R1516 AVDD.n1898 AVDD.n1897 2.18502
R1517 AVDD.n1893 AVDD.n1892 2.18502
R1518 AVDD.n1888 AVDD.n1887 2.18502
R1519 AVDD.n1806 AVDD.n1805 2.18502
R1520 AVDD.n1801 AVDD.n1800 2.18502
R1521 AVDD.n1796 AVDD.n1795 2.18502
R1522 AVDD.n1855 AVDD.n1854 2.18502
R1523 AVDD.n1850 AVDD.n1849 2.18502
R1524 AVDD.n1845 AVDD.n1844 2.18502
R1525 AVDD.n1840 AVDD.n1839 2.18502
R1526 AVDD.n1825 AVDD.n1824 2.18502
R1527 AVDD.n1820 AVDD.n1819 2.18502
R1528 AVDD.n1815 AVDD.n1814 2.18502
R1529 AVDD.n1485 AVDD.n1484 2.18502
R1530 AVDD.n1482 AVDD.n1481 2.18502
R1531 AVDD.n1479 AVDD.n1478 2.18502
R1532 AVDD.n1476 AVDD.n1475 2.18502
R1533 AVDD.n1471 AVDD.n1470 2.18502
R1534 AVDD.n1466 AVDD.n1465 2.18502
R1535 AVDD.n1461 AVDD.n1460 2.18502
R1536 AVDD.n1522 AVDD.n1521 2.18502
R1537 AVDD.n1519 AVDD.n1518 2.18502
R1538 AVDD.n1516 AVDD.n1515 2.18502
R1539 AVDD.n1513 AVDD.n1512 2.18502
R1540 AVDD.n1508 AVDD.n1507 2.18502
R1541 AVDD.n1503 AVDD.n1502 2.18502
R1542 AVDD.n1498 AVDD.n1497 2.18502
R1543 AVDD.n917 AVDD.n916 2.1566
R1544 AVDD.n914 AVDD.n913 2.1566
R1545 AVDD.n911 AVDD.n910 2.1566
R1546 AVDD.n906 AVDD.n905 2.1566
R1547 AVDD.n903 AVDD.n902 2.1566
R1548 AVDD.n682 AVDD.n681 2.14594
R1549 AVDD.n679 AVDD.n678 2.14594
R1550 AVDD.n676 AVDD.n675 2.14594
R1551 AVDD.n671 AVDD.n670 2.14594
R1552 AVDD.n668 AVDD.n667 2.14594
R1553 AVDD.n1866 AVDD.n1828 2.0852
R1554 AVDD.n1698 AVDD.n1653 2.0852
R1555 AVDD.n1535 AVDD.n1534 2.0852
R1556 AVDD.n212 AVDD.n211 2.0852
R1557 AVDD.n1922 AVDD.n1920 1.73609
R1558 AVDD.n1875 AVDD.n1785 1.73609
R1559 AVDD.n1599 AVDD.n1598 1.73609
R1560 AVDD.n1560 AVDD.n1559 1.73609
R1561 AVDD.n1758 AVDD.n1757 1.73383
R1562 AVDD.n1760 AVDD.n1759 1.73383
R1563 AVDD.n1763 AVDD.n1762 1.73383
R1564 AVDD.n1767 AVDD.n1766 1.73383
R1565 AVDD.n1771 AVDD.n1770 1.73383
R1566 AVDD.n1776 AVDD.n1775 1.73383
R1567 AVDD.n1778 AVDD.n1777 1.73383
R1568 AVDD.n1781 AVDD.n1780 1.73383
R1569 AVDD.n1309 AVDD.n1294 1.73383
R1570 AVDD.n1307 AVDD.n1295 1.73383
R1571 AVDD.n1304 AVDD.n1297 1.73383
R1572 AVDD.n1298 AVDD.n24 1.73383
R1573 AVDD.n1973 AVDD.n25 1.73383
R1574 AVDD.n1968 AVDD.n28 1.73383
R1575 AVDD.n1966 AVDD.n29 1.73383
R1576 AVDD.n1963 AVDD.n31 1.73383
R1577 AVDD.n1310 AVDD.n1309 1.73383
R1578 AVDD.n1307 AVDD.n1306 1.73383
R1579 AVDD.n1305 AVDD.n1304 1.73383
R1580 AVDD.n1300 AVDD.n24 1.73383
R1581 AVDD.n1973 AVDD.n1972 1.73383
R1582 AVDD.n1969 AVDD.n1968 1.73383
R1583 AVDD.n1966 AVDD.n1965 1.73383
R1584 AVDD.n1964 AVDD.n1963 1.73383
R1585 AVDD.n435 AVDD.n398 1.73383
R1586 AVDD.n433 AVDD.n399 1.73383
R1587 AVDD.n430 AVDD.n401 1.73383
R1588 AVDD.n425 AVDD.n403 1.73383
R1589 AVDD.n422 AVDD.n404 1.73383
R1590 AVDD.n417 AVDD.n407 1.73383
R1591 AVDD.n415 AVDD.n408 1.73383
R1592 AVDD.n412 AVDD.n410 1.73383
R1593 AVDD.n436 AVDD.n435 1.73383
R1594 AVDD.n433 AVDD.n432 1.73383
R1595 AVDD.n431 AVDD.n430 1.73383
R1596 AVDD.n426 AVDD.n425 1.73383
R1597 AVDD.n422 AVDD.n421 1.73383
R1598 AVDD.n418 AVDD.n417 1.73383
R1599 AVDD.n415 AVDD.n414 1.73383
R1600 AVDD.n413 AVDD.n412 1.73383
R1601 AVDD.n395 AVDD.n394 1.73383
R1602 AVDD.n392 AVDD.n391 1.73383
R1603 AVDD.n390 AVDD.n389 1.73383
R1604 AVDD.n385 AVDD.n384 1.73383
R1605 AVDD.n381 AVDD.n380 1.73383
R1606 AVDD.n377 AVDD.n376 1.73383
R1607 AVDD.n374 AVDD.n373 1.73383
R1608 AVDD.n372 AVDD.n371 1.73383
R1609 AVDD.n544 AVDD.n543 1.73383
R1610 AVDD.n541 AVDD.n540 1.73383
R1611 AVDD.n539 AVDD.n538 1.73383
R1612 AVDD.n534 AVDD.n533 1.73383
R1613 AVDD.n530 AVDD.n529 1.73383
R1614 AVDD.n526 AVDD.n525 1.73383
R1615 AVDD.n523 AVDD.n522 1.73383
R1616 AVDD.n521 AVDD.n520 1.73383
R1617 AVDD.n308 AVDD.n307 1.73383
R1618 AVDD.n305 AVDD.n304 1.73383
R1619 AVDD.n303 AVDD.n302 1.73383
R1620 AVDD.n298 AVDD.n82 1.73383
R1621 AVDD.n1440 AVDD.n1439 1.73383
R1622 AVDD.n1445 AVDD.n1444 1.73383
R1623 AVDD.n1447 AVDD.n1446 1.73383
R1624 AVDD.n1450 AVDD.n1449 1.73383
R1625 AVDD.n1324 AVDD.n1323 1.73383
R1626 AVDD.n1328 AVDD.n1327 1.73383
R1627 AVDD.n1330 AVDD.n1329 1.73383
R1628 AVDD.n1336 AVDD.n1335 1.73383
R1629 AVDD.n1338 AVDD.n1337 1.73383
R1630 AVDD.n1343 AVDD.n1342 1.73383
R1631 AVDD.n1347 AVDD.n1346 1.73383
R1632 AVDD.n1349 AVDD.n1348 1.73383
R1633 AVDD.n1325 AVDD.n1324 1.73383
R1634 AVDD.n1327 AVDD.n1326 1.73383
R1635 AVDD.n1331 AVDD.n1330 1.73383
R1636 AVDD.n1335 AVDD.n1334 1.73383
R1637 AVDD.n1339 AVDD.n1338 1.73383
R1638 AVDD.n1344 AVDD.n1343 1.73383
R1639 AVDD.n1346 AVDD.n1345 1.73383
R1640 AVDD.n1350 AVDD.n1349 1.73383
R1641 AVDD.n339 AVDD.n324 1.73383
R1642 AVDD.n337 AVDD.n325 1.73383
R1643 AVDD.n334 AVDD.n327 1.73383
R1644 AVDD.n328 AVDD.n93 1.73383
R1645 AVDD.n1431 AVDD.n94 1.73383
R1646 AVDD.n1426 AVDD.n97 1.73383
R1647 AVDD.n1424 AVDD.n98 1.73383
R1648 AVDD.n1421 AVDD.n100 1.73383
R1649 AVDD.n340 AVDD.n339 1.73383
R1650 AVDD.n337 AVDD.n336 1.73383
R1651 AVDD.n335 AVDD.n334 1.73383
R1652 AVDD.n330 AVDD.n93 1.73383
R1653 AVDD.n1431 AVDD.n1430 1.73383
R1654 AVDD.n1427 AVDD.n1426 1.73383
R1655 AVDD.n1424 AVDD.n1423 1.73383
R1656 AVDD.n1422 AVDD.n1421 1.73383
R1657 AVDD.n567 AVDD.n566 1.73383
R1658 AVDD.n571 AVDD.n570 1.73383
R1659 AVDD.n573 AVDD.n572 1.73383
R1660 AVDD.n579 AVDD.n578 1.73383
R1661 AVDD.n581 AVDD.n580 1.73383
R1662 AVDD.n586 AVDD.n585 1.73383
R1663 AVDD.n590 AVDD.n589 1.73383
R1664 AVDD.n592 AVDD.n591 1.73383
R1665 AVDD.n602 AVDD.n601 1.73383
R1666 AVDD.n606 AVDD.n605 1.73383
R1667 AVDD.n608 AVDD.n607 1.73383
R1668 AVDD.n611 AVDD.n114 1.73383
R1669 AVDD.n1390 AVDD.n115 1.73383
R1670 AVDD.n1385 AVDD.n616 1.73383
R1671 AVDD.n1383 AVDD.n617 1.73383
R1672 AVDD.n1380 AVDD.n619 1.73383
R1673 AVDD.n568 AVDD.n567 1.73383
R1674 AVDD.n570 AVDD.n569 1.73383
R1675 AVDD.n574 AVDD.n573 1.73383
R1676 AVDD.n578 AVDD.n577 1.73383
R1677 AVDD.n582 AVDD.n581 1.73383
R1678 AVDD.n587 AVDD.n586 1.73383
R1679 AVDD.n589 AVDD.n588 1.73383
R1680 AVDD.n593 AVDD.n592 1.73383
R1681 AVDD.n603 AVDD.n602 1.73383
R1682 AVDD.n605 AVDD.n604 1.73383
R1683 AVDD.n609 AVDD.n608 1.73383
R1684 AVDD.n614 AVDD.n114 1.73383
R1685 AVDD.n1390 AVDD.n1389 1.73383
R1686 AVDD.n1386 AVDD.n1385 1.73383
R1687 AVDD.n1383 AVDD.n1382 1.73383
R1688 AVDD.n1381 AVDD.n1380 1.73383
R1689 AVDD.n474 AVDD.n473 1.73383
R1690 AVDD.n478 AVDD.n477 1.73383
R1691 AVDD.n480 AVDD.n479 1.73383
R1692 AVDD.n486 AVDD.n485 1.73383
R1693 AVDD.n488 AVDD.n487 1.73383
R1694 AVDD.n493 AVDD.n492 1.73383
R1695 AVDD.n497 AVDD.n496 1.73383
R1696 AVDD.n499 AVDD.n498 1.73383
R1697 AVDD.n475 AVDD.n474 1.73383
R1698 AVDD.n477 AVDD.n476 1.73383
R1699 AVDD.n481 AVDD.n480 1.73383
R1700 AVDD.n485 AVDD.n484 1.73383
R1701 AVDD.n489 AVDD.n488 1.73383
R1702 AVDD.n494 AVDD.n493 1.73383
R1703 AVDD.n496 AVDD.n495 1.73383
R1704 AVDD.n500 AVDD.n499 1.73383
R1705 AVDD.n1145 AVDD.n1144 1.73383
R1706 AVDD.n1991 AVDD.n1990 1.73383
R1707 AVDD.n1988 AVDD.n1987 1.73383
R1708 AVDD.n1986 AVDD.n1985 1.73383
R1709 AVDD.n1981 AVDD.n1980 1.73383
R1710 AVDD.n852 AVDD.n851 1.73383
R1711 AVDD.n856 AVDD.n855 1.73383
R1712 AVDD.n861 AVDD.n860 1.73383
R1713 AVDD.n778 AVDD.n730 1.73383
R1714 AVDD.n776 AVDD.n731 1.73383
R1715 AVDD.n773 AVDD.n733 1.73383
R1716 AVDD.n768 AVDD.n735 1.73383
R1717 AVDD.n765 AVDD.n736 1.73383
R1718 AVDD.n760 AVDD.n739 1.73383
R1719 AVDD.n758 AVDD.n740 1.73383
R1720 AVDD.n755 AVDD.n742 1.73383
R1721 AVDD.n779 AVDD.n778 1.73383
R1722 AVDD.n776 AVDD.n775 1.73383
R1723 AVDD.n774 AVDD.n773 1.73383
R1724 AVDD.n769 AVDD.n768 1.73383
R1725 AVDD.n765 AVDD.n764 1.73383
R1726 AVDD.n761 AVDD.n760 1.73383
R1727 AVDD.n758 AVDD.n757 1.73383
R1728 AVDD.n756 AVDD.n755 1.73383
R1729 AVDD.n794 AVDD.n793 1.73383
R1730 AVDD.n798 AVDD.n797 1.73383
R1731 AVDD.n800 AVDD.n799 1.73383
R1732 AVDD.n806 AVDD.n805 1.73383
R1733 AVDD.n808 AVDD.n807 1.73383
R1734 AVDD.n813 AVDD.n812 1.73383
R1735 AVDD.n817 AVDD.n816 1.73383
R1736 AVDD.n819 AVDD.n818 1.73383
R1737 AVDD.n795 AVDD.n794 1.73383
R1738 AVDD.n797 AVDD.n796 1.73383
R1739 AVDD.n801 AVDD.n800 1.73383
R1740 AVDD.n805 AVDD.n804 1.73383
R1741 AVDD.n809 AVDD.n808 1.73383
R1742 AVDD.n814 AVDD.n813 1.73383
R1743 AVDD.n816 AVDD.n815 1.73383
R1744 AVDD.n820 AVDD.n819 1.73383
R1745 AVDD.n1001 AVDD.n1000 1.73383
R1746 AVDD.n1003 AVDD.n1002 1.73383
R1747 AVDD.n1006 AVDD.n1005 1.73383
R1748 AVDD.n1010 AVDD.n1009 1.73383
R1749 AVDD.n1014 AVDD.n1013 1.73383
R1750 AVDD.n1019 AVDD.n1018 1.73383
R1751 AVDD.n1021 AVDD.n1020 1.73383
R1752 AVDD.n1024 AVDD.n1023 1.73383
R1753 AVDD.n872 AVDD.n871 1.73383
R1754 AVDD.n874 AVDD.n873 1.73383
R1755 AVDD.n879 AVDD.n878 1.73383
R1756 AVDD.n885 AVDD.n695 1.73383
R1757 AVDD.n886 AVDD.n698 1.73383
R1758 AVDD.n722 AVDD.n721 1.73383
R1759 AVDD.n708 AVDD.n706 1.73383
R1760 AVDD.n714 AVDD.n713 1.73383
R1761 AVDD.n865 AVDD.n864 1.73383
R1762 AVDD.n883 AVDD.n882 1.73383
R1763 AVDD.n893 AVDD.n892 1.73383
R1764 AVDD.n891 AVDD.n890 1.73383
R1765 AVDD.n720 AVDD.n719 1.73383
R1766 AVDD.n718 AVDD.n717 1.73383
R1767 AVDD.n1140 AVDD.n1139 1.73383
R1768 AVDD.n1142 AVDD.n1141 1.73383
R1769 AVDD.n1174 AVDD.n1173 1.73383
R1770 AVDD.n1178 AVDD.n1177 1.73383
R1771 AVDD.n1180 AVDD.n1179 1.73383
R1772 AVDD.n1186 AVDD.n1185 1.73383
R1773 AVDD.n1188 AVDD.n1187 1.73383
R1774 AVDD.n1193 AVDD.n1192 1.73383
R1775 AVDD.n1197 AVDD.n1196 1.73383
R1776 AVDD.n1199 AVDD.n1198 1.73383
R1777 AVDD.n1175 AVDD.n1174 1.73383
R1778 AVDD.n1177 AVDD.n1176 1.73383
R1779 AVDD.n1181 AVDD.n1180 1.73383
R1780 AVDD.n1185 AVDD.n1184 1.73383
R1781 AVDD.n1189 AVDD.n1188 1.73383
R1782 AVDD.n1194 AVDD.n1193 1.73383
R1783 AVDD.n1196 AVDD.n1195 1.73383
R1784 AVDD.n1200 AVDD.n1199 1.73383
R1785 AVDD.n1290 AVDD.n621 1.73383
R1786 AVDD.n1288 AVDD.n622 1.73383
R1787 AVDD.n1285 AVDD.n624 1.73383
R1788 AVDD.n1280 AVDD.n626 1.73383
R1789 AVDD.n1277 AVDD.n627 1.73383
R1790 AVDD.n1272 AVDD.n630 1.73383
R1791 AVDD.n1270 AVDD.n631 1.73383
R1792 AVDD.n1267 AVDD.n633 1.73383
R1793 AVDD.n1254 AVDD.n638 1.73383
R1794 AVDD.n1252 AVDD.n639 1.73383
R1795 AVDD.n1249 AVDD.n641 1.73383
R1796 AVDD.n1244 AVDD.n643 1.73383
R1797 AVDD.n1241 AVDD.n645 1.73383
R1798 AVDD.n1236 AVDD.n648 1.73383
R1799 AVDD.n1234 AVDD.n649 1.73383
R1800 AVDD.n1231 AVDD.n651 1.73383
R1801 AVDD.n1291 AVDD.n1290 1.73383
R1802 AVDD.n1288 AVDD.n1287 1.73383
R1803 AVDD.n1286 AVDD.n1285 1.73383
R1804 AVDD.n1281 AVDD.n1280 1.73383
R1805 AVDD.n1277 AVDD.n1276 1.73383
R1806 AVDD.n1273 AVDD.n1272 1.73383
R1807 AVDD.n1270 AVDD.n1269 1.73383
R1808 AVDD.n1268 AVDD.n1267 1.73383
R1809 AVDD.n1255 AVDD.n1254 1.73383
R1810 AVDD.n1252 AVDD.n1251 1.73383
R1811 AVDD.n1250 AVDD.n1249 1.73383
R1812 AVDD.n1245 AVDD.n1244 1.73383
R1813 AVDD.n1241 AVDD.n1240 1.73383
R1814 AVDD.n1237 AVDD.n1236 1.73383
R1815 AVDD.n1234 AVDD.n1233 1.73383
R1816 AVDD.n1232 AVDD.n1231 1.73383
R1817 AVDD.n1633 AVDD.n1632 1.73383
R1818 AVDD.n1631 AVDD.n1630 1.73383
R1819 AVDD.n1628 AVDD.n1627 1.73383
R1820 AVDD.n1624 AVDD.n1623 1.73383
R1821 AVDD.n1620 AVDD.n1619 1.73383
R1822 AVDD.n1616 AVDD.n1615 1.73383
R1823 AVDD.n1613 AVDD.n1612 1.73383
R1824 AVDD.n1934 AVDD.n1933 1.73383
R1825 AVDD.n174 AVDD.n173 1.73383
R1826 AVDD.n172 AVDD.n171 1.73383
R1827 AVDD.n169 AVDD.n168 1.73383
R1828 AVDD.n165 AVDD.n164 1.73383
R1829 AVDD.n161 AVDD.n160 1.73383
R1830 AVDD.n157 AVDD.n156 1.73383
R1831 AVDD.n154 AVDD.n153 1.73383
R1832 AVDD.n1603 AVDD.n1602 1.73383
R1833 AVDD.n1748 AVDD.n1634 1.69136
R1834 AVDD.n1756 AVDD.n1755 1.69136
R1835 AVDD.n289 AVDD.n175 1.69136
R1836 AVDD.n295 AVDD.n294 1.69136
R1837 AVDD.n1747 AVDD.n1746 1.65018
R1838 AVDD.n1669 AVDD.n1665 1.65018
R1839 AVDD.n259 AVDD.n143 1.65018
R1840 AVDD.n230 AVDD.n229 1.65018
R1841 AVDD.n1605 AVDD.t432 1.60217
R1842 AVDD.n2022 AVDD.t954 1.60217
R1843 AVDD.n2019 AVDD.t855 1.60217
R1844 AVDD.n2 AVDD.t924 1.60217
R1845 AVDD.n1354 AVDD.t1106 1.60217
R1846 AVDD.n1356 AVDD.t350 1.60217
R1847 AVDD.n1605 AVDD.t1188 1.60217
R1848 AVDD.n2022 AVDD.t416 1.60217
R1849 AVDD.n2019 AVDD.t321 1.60217
R1850 AVDD.n2 AVDD.t392 1.60217
R1851 AVDD.n1354 AVDD.t588 1.60217
R1852 AVDD.n1356 AVDD.t1084 1.60217
R1853 AVDD.n1358 AVDD.t982 1.60217
R1854 AVDD.n1360 AVDD.t208 1.60217
R1855 AVDD.n1363 AVDD.t71 1.60217
R1856 AVDD.n1366 AVDD.t212 1.60217
R1857 AVDD.n1369 AVDD.t73 1.60217
R1858 AVDD.n1371 AVDD.t677 1.60217
R1859 AVDD.n1358 AVDD.t442 1.60217
R1860 AVDD.n1360 AVDD.t960 1.60217
R1861 AVDD.n1363 AVDD.t867 1.60217
R1862 AVDD.n1366 AVDD.t222 1.60217
R1863 AVDD.n1369 AVDD.t115 1.60217
R1864 AVDD.n1371 AVDD.t695 1.60217
R1865 AVDD.n1376 AVDD.t681 1.60217
R1866 AVDD.n1374 AVDD.t1178 1.60217
R1867 AVDD.n10 AVDD.t1060 1.60217
R1868 AVDD.n2013 AVDD.t1066 1.60217
R1869 AVDD.n2010 AVDD.t760 1.60217
R1870 AVDD.n2008 AVDD.t849 1.60217
R1871 AVDD.n1376 AVDD.t703 1.60217
R1872 AVDD.n1374 AVDD.t1192 1.60217
R1873 AVDD.n10 AVDD.t1070 1.60217
R1874 AVDD.n2013 AVDD.t1090 1.60217
R1875 AVDD.n2010 AVDD.t262 1.60217
R1876 AVDD.n2008 AVDD.t315 1.60217
R1877 AVDD.n2006 AVDD.t1226 1.60217
R1878 AVDD.n2004 AVDD.t669 1.60217
R1879 AVDD.n2001 AVDD.t794 1.60217
R1880 AVDD.n1999 AVDD.t782 1.60217
R1881 AVDD.n1996 AVDD.t890 1.60217
R1882 AVDD.n1994 AVDD.t371 1.60217
R1883 AVDD.n2006 AVDD.t726 1.60217
R1884 AVDD.n2004 AVDD.t129 1.60217
R1885 AVDD.n2001 AVDD.t267 1.60217
R1886 AVDD.n1999 AVDD.t248 1.60217
R1887 AVDD.n1996 AVDD.t354 1.60217
R1888 AVDD.n1994 AVDD.t1120 1.60217
R1889 AVDD.n1937 AVDD.t47 1.60217
R1890 AVDD.n1939 AVDD.t584 1.60217
R1891 AVDD.n1942 AVDD.t452 1.60217
R1892 AVDD.n1948 AVDD.t551 1.60217
R1893 AVDD.n1945 AVDD.t752 1.60217
R1894 AVDD.n33 AVDD.t1236 1.60217
R1895 AVDD.n1937 AVDD.t169 1.60217
R1896 AVDD.n1939 AVDD.t691 1.60217
R1897 AVDD.n1942 AVDD.t578 1.60217
R1898 AVDD.n1948 AVDD.t651 1.60217
R1899 AVDD.n1945 AVDD.t863 1.60217
R1900 AVDD.n33 AVDD.t49 1.60217
R1901 AVDD.n1959 AVDD.t606 1.60217
R1902 AVDD.n1957 AVDD.t1100 1.60217
R1903 AVDD.n1954 AVDD.t1000 1.60217
R1904 AVDD.n34 AVDD.t882 1.60217
R1905 AVDD.n1261 AVDD.t774 1.60217
R1906 AVDD.n1959 AVDD.t720 1.60217
R1907 AVDD.n1957 AVDD.t1206 1.60217
R1908 AVDD.n1954 AVDD.t1096 1.60217
R1909 AVDD.n34 AVDD.t458 1.60217
R1910 AVDD.n1261 AVDD.t358 1.60217
R1911 AVDD.n1225 AVDD.t626 1.60217
R1912 AVDD.n1222 AVDD.t515 1.60217
R1913 AVDD.n654 AVDD.t521 1.60217
R1914 AVDD.n749 AVDD.t1196 1.60217
R1915 AVDD.n1211 AVDD.t1130 1.60217
R1916 AVDD.n1208 AVDD.t1014 1.60217
R1917 AVDD.n1206 AVDD.t936 1.60217
R1918 AVDD.n653 AVDD.t833 1.60217
R1919 AVDD.n56 AVDD.t63 1.60217
R1920 AVDD.n1156 AVDD.t596 1.60217
R1921 AVDD.n1159 AVDD.t487 1.60217
R1922 AVDD.n1216 AVDD.t564 1.60217
R1923 AVDD.n1213 AVDD.t776 1.60217
R1924 AVDD.n468 AVDD.t1256 1.60217
R1925 AVDD.n356 AVDD.t101 1.60217
R1926 AVDD.n551 AVDD.t68 1.60217
R1927 AVDD.n548 AVDD.t203 1.60217
R1928 AVDD.n546 AVDD.t980 1.60217
R1929 AVDD.n561 AVDD.t1094 1.60217
R1930 AVDD.n558 AVDD.t998 1.60217
R1931 AVDD.n462 AVDD.t1004 1.60217
R1932 AVDD.n465 AVDD.t636 1.60217
R1933 AVDD.n125 AVDD.t198 1.60217
R1934 AVDD.n440 AVDD.t57 1.60217
R1935 AVDD.n443 AVDD.t75 1.60217
R1936 AVDD.n446 AVDD.t547 1.60217
R1937 AVDD.n448 AVDD.t604 1.60217
R1938 AVDD.n125 AVDD.t930 1.60217
R1939 AVDD.n440 AVDD.t825 1.60217
R1940 AVDD.n443 AVDD.t843 1.60217
R1941 AVDD.n446 AVDD.t831 1.60217
R1942 AVDD.n448 AVDD.t163 1.60217
R1943 AVDD.n503 AVDD.t1002 1.60217
R1944 AVDD.n505 AVDD.t420 1.60217
R1945 AVDD.n508 AVDD.t545 1.60217
R1946 AVDD.n511 AVDD.t529 1.60217
R1947 AVDD.n514 AVDD.t634 1.60217
R1948 AVDD.n516 AVDD.t127 1.60217
R1949 AVDD.n503 AVDD.t582 1.60217
R1950 AVDD.n505 AVDD.t1258 1.60217
R1951 AVDD.n508 AVDD.t109 1.60217
R1952 AVDD.n511 AVDD.t80 1.60217
R1953 AVDD.n514 AVDD.t214 1.60217
R1954 AVDD.n516 AVDD.t990 1.60217
R1955 AVDD.n1396 AVDD.t210 1.60217
R1956 AVDD.n1398 AVDD.t730 1.60217
R1957 AVDD.n1401 AVDD.t608 1.60217
R1958 AVDD.n1406 AVDD.t685 1.60217
R1959 AVDD.n1403 AVDD.t894 1.60217
R1960 AVDD.n102 AVDD.t96 1.60217
R1961 AVDD.n1396 AVDD.t1050 1.60217
R1962 AVDD.n1398 AVDD.t301 1.60217
R1963 AVDD.n1401 AVDD.t167 1.60217
R1964 AVDD.n1406 AVDD.t271 1.60217
R1965 AVDD.n1403 AVDD.t440 1.60217
R1966 AVDD.n102 AVDD.t958 1.60217
R1967 AVDD.n1417 AVDD.t754 1.60217
R1968 AVDD.n1415 AVDD.t1238 1.60217
R1969 AVDD.n1412 AVDD.t1144 1.60217
R1970 AVDD.n103 AVDD.t499 1.60217
R1971 AVDD.n124 AVDD.t390 1.60217
R1972 AVDD.n1417 AVDD.t319 1.60217
R1973 AVDD.n1415 AVDD.t837 1.60217
R1974 AVDD.n1412 AVDD.t722 1.60217
R1975 AVDD.n103 AVDD.t1220 1.60217
R1976 AVDD.n124 AVDD.t1116 1.60217
R1977 AVDD.n345 AVDD.t823 1.60217
R1978 AVDD.n348 AVDD.t711 1.60217
R1979 AVDD.n351 AVDD.t125 1.60217
R1980 AVDD.n354 AVDD.t1272 1.60217
R1981 AVDD.n310 AVDD.t1038 1.60217
R1982 AVDD.n312 AVDD.t297 1.60217
R1983 AVDD.n315 AVDD.t159 1.60217
R1984 AVDD.n318 AVDD.t260 1.60217
R1985 AVDD.n321 AVDD.t428 1.60217
R1986 AVDD.n694 AVDD.t1080 1.60217
R1987 AVDD.n938 AVDD.t659 1.60217
R1988 AVDD.n1050 AVDD.t784 1.60217
R1989 AVDD.n928 AVDD.t191 1.60217
R1990 AVDD.n1122 AVDD.t946 1.60217
R1991 AVDD.n1119 AVDD.t132 1.60217
R1992 AVDD.n693 AVDD.t679 1.60217
R1993 AVDD.n746 AVDD.t313 1.60217
R1994 AVDD.n659 AVDD.t414 1.60217
R1995 AVDD.n1152 AVDD.t406 1.60217
R1996 AVDD.n1149 AVDD.t517 1.60217
R1997 AVDD.n1147 AVDD.t1262 1.60217
R1998 AVDD.n635 AVDD.t566 1.60217
R1999 AVDD.n824 AVDD.t438 1.60217
R2000 AVDD.n827 AVDD.t450 1.60217
R2001 AVDD.n830 AVDD.t1018 1.60217
R2002 AVDD.n832 AVDD.t448 1.60217
R2003 AVDD.n635 AVDD.t144 1.60217
R2004 AVDD.n824 AVDD.t17 1.60217
R2005 AVDD.n827 AVDD.t42 1.60217
R2006 AVDD.n830 AVDD.t701 1.60217
R2007 AVDD.n832 AVDD.t574 1.60217
R2008 AVDD.n834 AVDD.t878 1.60217
R2009 AVDD.n836 AVDD.t303 1.60217
R2010 AVDD.n839 AVDD.t402 1.60217
R2011 AVDD.n841 AVDD.t386 1.60217
R2012 AVDD.n844 AVDD.t497 1.60217
R2013 AVDD.n834 AVDD.t978 1.60217
R2014 AVDD.n836 AVDD.t397 1.60217
R2015 AVDD.n839 AVDD.t513 1.60217
R2016 AVDD.n841 AVDD.t493 1.60217
R2017 AVDD.n844 AVDD.t614 1.60217
R2018 AVDD.n663 AVDD.t984 1.60217
R2019 AVDD.n685 AVDD.t182 1.60217
R2020 AVDD.n1097 AVDD.t724 1.60217
R2021 AVDD.n941 AVDD.t1142 1.60217
R2022 AVDD.n945 AVDD.t707 1.60217
R2023 AVDD.n918 AVDD.t817 1.60217
R2024 AVDD.n1026 AVDD.t246 1.60217
R2025 AVDD.n1906 AVDD.n1905 1.60175
R2026 AVDD.n1562 AVDD.n1561 1.60175
R2027 AVDD.n1129 AVDD.n1127 1.57603
R2028 AVDD.n955 AVDD.n953 1.57603
R2029 AVDD.n1912 AVDD.n46 1.5005
R2030 AVDD.n1883 AVDD.n1882 1.5005
R2031 AVDD.n1885 AVDD.n1884 1.5005
R2032 AVDD.n1930 AVDD.n1929 1.5005
R2033 AVDD.n1866 AVDD.n1865 1.5005
R2034 AVDD.n1705 AVDD.n1704 1.5005
R2035 AVDD.n1707 AVDD.n1706 1.5005
R2036 AVDD.n1755 AVDD.n1754 1.5005
R2037 AVDD.n1698 AVDD.n1697 1.5005
R2038 AVDD.n1730 AVDD.n63 1.5005
R2039 AVDD.n1536 AVDD.n1535 1.5005
R2040 AVDD.n1588 AVDD.n1587 1.5005
R2041 AVDD.n1551 AVDD.n1454 1.5005
R2042 AVDD.n1575 AVDD.n1574 1.5005
R2043 AVDD.n1590 AVDD.n1589 1.5005
R2044 AVDD.n233 AVDD.n176 1.5005
R2045 AVDD.n255 AVDD.n254 1.5005
R2046 AVDD.n290 AVDD.n289 1.5005
R2047 AVDD.n213 AVDD.n212 1.5005
R2048 AVDD.n288 AVDD.n287 1.5005
R2049 AVDD.n1603 AVDD.t1008 1.4705
R2050 AVDD.t139 AVDD.n1603 1.4705
R2051 AVDD.n153 AVDD.t1264 1.4705
R2052 AVDD.n153 AVDD.t1008 1.4705
R2053 AVDD.t422 AVDD.n157 1.4705
R2054 AVDD.n157 AVDD.t1264 1.4705
R2055 AVDD.n160 AVDD.t671 1.4705
R2056 AVDD.n160 AVDD.t384 1.4705
R2057 AVDD.t1076 AVDD.n165 1.4705
R2058 AVDD.n165 AVDD.t671 1.4705
R2059 AVDD.n168 AVDD.t112 1.4705
R2060 AVDD.n168 AVDD.t1108 1.4705
R2061 AVDD.t653 AVDD.n172 1.4705
R2062 AVDD.n172 AVDD.t112 1.4705
R2063 AVDD.n173 AVDD.t934 1.4705
R2064 AVDD.n173 AVDD.t653 1.4705
R2065 AVDD.n1934 AVDD.t948 1.4705
R2066 AVDD.t1208 AVDD.n1934 1.4705
R2067 AVDD.n1612 AVDD.t54 1.4705
R2068 AVDD.n1612 AVDD.t948 1.4705
R2069 AVDD.t1064 AVDD.n1616 1.4705
R2070 AVDD.n1616 AVDD.t54 1.4705
R2071 AVDD.n1619 AVDD.t713 1.4705
R2072 AVDD.n1619 AVDD.t1136 1.4705
R2073 AVDD.t418 AVDD.n1624 1.4705
R2074 AVDD.n1624 AVDD.t713 1.4705
R2075 AVDD.n1627 AVDD.t269 1.4705
R2076 AVDD.n1627 AVDD.t287 1.4705
R2077 AVDD.t643 AVDD.n1631 1.4705
R2078 AVDD.n1631 AVDD.t269 1.4705
R2079 AVDD.n1632 AVDD.t1168 1.4705
R2080 AVDD.n1632 AVDD.t643 1.4705
R2081 AVDD.t285 AVDD.n1232 1.4705
R2082 AVDD.n1232 AVDD.t665 1.4705
R2083 AVDD.n1233 AVDD.t966 1.4705
R2084 AVDD.n1233 AVDD.t285 1.4705
R2085 AVDD.t904 AVDD.n1237 1.4705
R2086 AVDD.n1237 AVDD.t966 1.4705
R2087 AVDD.n1240 AVDD.t906 1.4705
R2088 AVDD.n1240 AVDD.t527 1.4705
R2089 AVDD.t501 AVDD.n1245 1.4705
R2090 AVDD.n1245 AVDD.t906 1.4705
R2091 AVDD.t472 AVDD.n1250 1.4705
R2092 AVDD.n1250 AVDD.t91 1.4705
R2093 AVDD.n1251 AVDD.t748 1.4705
R2094 AVDD.n1251 AVDD.t472 1.4705
R2095 AVDD.t1098 AVDD.n1255 1.4705
R2096 AVDD.n1255 AVDD.t748 1.4705
R2097 AVDD.t1068 AVDD.n1268 1.4705
R2098 AVDD.n1268 AVDD.t1158 1.4705
R2099 AVDD.n1269 AVDD.t495 1.4705
R2100 AVDD.n1269 AVDD.t1068 1.4705
R2101 AVDD.t426 AVDD.n1273 1.4705
R2102 AVDD.n1273 AVDD.t495 1.4705
R2103 AVDD.n1276 AVDD.t99 1.4705
R2104 AVDD.n1276 AVDD.t1016 1.4705
R2105 AVDD.t6 AVDD.n1281 1.4705
R2106 AVDD.n1281 AVDD.t99 1.4705
R2107 AVDD.t1036 AVDD.n1286 1.4705
R2108 AVDD.n1286 AVDD.t594 1.4705
R2109 AVDD.n1287 AVDD.t1126 1.4705
R2110 AVDD.n1287 AVDD.t1036 1.4705
R2111 AVDD.t1210 AVDD.n1291 1.4705
R2112 AVDD.n1291 AVDD.t1126 1.4705
R2113 AVDD.n651 AVDD.t289 1.4705
R2114 AVDD.t673 AVDD.n651 1.4705
R2115 AVDD.n649 AVDD.t972 1.4705
R2116 AVDD.t289 AVDD.n649 1.4705
R2117 AVDD.n648 AVDD.t910 1.4705
R2118 AVDD.t972 AVDD.n648 1.4705
R2119 AVDD.n645 AVDD.t912 1.4705
R2120 AVDD.t533 AVDD.n645 1.4705
R2121 AVDD.n643 AVDD.t509 1.4705
R2122 AVDD.t912 AVDD.n643 1.4705
R2123 AVDD.n641 AVDD.t485 1.4705
R2124 AVDD.t103 AVDD.n641 1.4705
R2125 AVDD.n639 AVDD.t756 1.4705
R2126 AVDD.t485 AVDD.n639 1.4705
R2127 AVDD.n638 AVDD.t1104 1.4705
R2128 AVDD.t756 AVDD.n638 1.4705
R2129 AVDD.n633 AVDD.t1082 1.4705
R2130 AVDD.t1166 AVDD.n633 1.4705
R2131 AVDD.n631 AVDD.t503 1.4705
R2132 AVDD.t1082 AVDD.n631 1.4705
R2133 AVDD.n630 AVDD.t430 1.4705
R2134 AVDD.t503 AVDD.n630 1.4705
R2135 AVDD.n627 AVDD.t107 1.4705
R2136 AVDD.t1020 AVDD.n627 1.4705
R2137 AVDD.n626 AVDD.t11 1.4705
R2138 AVDD.t107 AVDD.n626 1.4705
R2139 AVDD.n624 AVDD.t1046 1.4705
R2140 AVDD.t600 AVDD.n624 1.4705
R2141 AVDD.n622 AVDD.t1134 1.4705
R2142 AVDD.t1046 AVDD.n622 1.4705
R2143 AVDD.n621 AVDD.t1216 1.4705
R2144 AVDD.t1134 AVDD.n621 1.4705
R2145 AVDD.n1200 AVDD.t766 1.4705
R2146 AVDD.t715 AVDD.n1200 1.4705
R2147 AVDD.n1195 AVDD.t1170 1.4705
R2148 AVDD.n1195 AVDD.t766 1.4705
R2149 AVDD.n1194 AVDD.t900 1.4705
R2150 AVDD.t1170 AVDD.n1194 1.4705
R2151 AVDD.n1189 AVDD.t187 1.4705
R2152 AVDD.t620 AVDD.n1189 1.4705
R2153 AVDD.n1184 AVDD.t239 1.4705
R2154 AVDD.n1184 AVDD.t187 1.4705
R2155 AVDD.n1181 AVDD.t37 1.4705
R2156 AVDD.t489 AVDD.n1181 1.4705
R2157 AVDD.n1176 AVDD.t628 1.4705
R2158 AVDD.n1176 AVDD.t37 1.4705
R2159 AVDD.n1175 AVDD.t206 1.4705
R2160 AVDD.t628 AVDD.n1175 1.4705
R2161 AVDD.n1781 AVDD.t869 1.4705
R2162 AVDD.t819 AVDD.n1781 1.4705
R2163 AVDD.n1777 AVDD.t1248 1.4705
R2164 AVDD.n1777 AVDD.t869 1.4705
R2165 AVDD.n1776 AVDD.t996 1.4705
R2166 AVDD.t1248 AVDD.n1776 1.4705
R2167 AVDD.n1771 AVDD.t305 1.4705
R2168 AVDD.t732 AVDD.n1771 1.4705
R2169 AVDD.n1766 AVDD.t343 1.4705
R2170 AVDD.n1766 AVDD.t305 1.4705
R2171 AVDD.n1763 AVDD.t146 1.4705
R2172 AVDD.t586 AVDD.n1763 1.4705
R2173 AVDD.n1759 AVDD.t738 1.4705
R2174 AVDD.n1759 AVDD.t146 1.4705
R2175 AVDD.n1758 AVDD.t311 1.4705
R2176 AVDD.t738 AVDD.n1758 1.4705
R2177 AVDD.n1861 AVDD.t1652 1.4705
R2178 AVDD.n1861 AVDD.t1584 1.4705
R2179 AVDD.n1862 AVDD.t1374 1.4705
R2180 AVDD.n1862 AVDD.t1493 1.4705
R2181 AVDD.n1829 AVDD.t1421 1.4705
R2182 AVDD.n1829 AVDD.t1395 1.4705
R2183 AVDD.n1830 AVDD.t1665 1.4705
R2184 AVDD.n1830 AVDD.t1657 1.4705
R2185 AVDD.n1921 AVDD.t1420 1.4705
R2186 AVDD.n1921 AVDD.t1642 1.4705
R2187 AVDD.n1923 AVDD.t1411 1.4705
R2188 AVDD.n1923 AVDD.t1478 1.4705
R2189 AVDD.n1925 AVDD.t1467 1.4705
R2190 AVDD.n1925 AVDD.t1687 1.4705
R2191 AVDD.n1927 AVDD.t1673 1.4705
R2192 AVDD.n1927 AVDD.t1580 1.4705
R2193 AVDD.n52 AVDD.t1433 1.4705
R2194 AVDD.n52 AVDD.t1491 1.4705
R2195 AVDD.n50 AVDD.t1402 1.4705
R2196 AVDD.n50 AVDD.t1446 1.4705
R2197 AVDD.n48 AVDD.t1297 1.4705
R2198 AVDD.n48 AVDD.t1294 1.4705
R2199 AVDD.n47 AVDD.t1386 1.4705
R2200 AVDD.n47 AVDD.t1678 1.4705
R2201 AVDD.n1902 AVDD.t1409 1.4705
R2202 AVDD.n1902 AVDD.t1430 1.4705
R2203 AVDD.n1897 AVDD.t1389 1.4705
R2204 AVDD.n1897 AVDD.t1470 1.4705
R2205 AVDD.n1892 AVDD.t1669 1.4705
R2206 AVDD.n1892 AVDD.t1655 1.4705
R2207 AVDD.n1887 AVDD.t1572 1.4705
R2208 AVDD.n1887 AVDD.t1439 1.4705
R2209 AVDD.n1805 AVDD.t1398 1.4705
R2210 AVDD.n1805 AVDD.t1443 1.4705
R2211 AVDD.n1800 AVDD.t1487 1.4705
R2212 AVDD.n1800 AVDD.t1301 1.4705
R2213 AVDD.n1795 AVDD.t1659 1.4705
R2214 AVDD.n1795 AVDD.t1577 1.4705
R2215 AVDD.n1793 AVDD.t1452 1.4705
R2216 AVDD.n1793 AVDD.t1643 1.4705
R2217 AVDD.n1874 AVDD.t1442 1.4705
R2218 AVDD.n1874 AVDD.t1449 1.4705
R2219 AVDD.n1876 AVDD.t1299 1.4705
R2220 AVDD.n1876 AVDD.t1564 1.4705
R2221 AVDD.n1878 AVDD.t1591 1.4705
R2222 AVDD.n1878 AVDD.t1396 1.4705
R2223 AVDD.n1880 AVDD.t1423 1.4705
R2224 AVDD.n1880 AVDD.t1482 1.4705
R2225 AVDD.n1872 AVDD.t1464 1.4705
R2226 AVDD.n1872 AVDD.t1570 1.4705
R2227 AVDD.n1870 AVDD.t1668 1.4705
R2228 AVDD.n1870 AVDD.t1681 1.4705
R2229 AVDD.n1868 AVDD.t1648 1.4705
R2230 AVDD.n1868 AVDD.t1644 1.4705
R2231 AVDD.n1867 AVDD.t1579 1.4705
R2232 AVDD.n1867 AVDD.t1385 1.4705
R2233 AVDD.n1854 AVDD.t1571 1.4705
R2234 AVDD.n1854 AVDD.t1419 1.4705
R2235 AVDD.n1849 AVDD.t1400 1.4705
R2236 AVDD.n1849 AVDD.t1388 1.4705
R2237 AVDD.n1844 AVDD.t1596 1.4705
R2238 AVDD.n1844 AVDD.t1286 1.4705
R2239 AVDD.n1839 AVDD.t1456 1.4705
R2240 AVDD.n1839 AVDD.t1435 1.4705
R2241 AVDD.n1824 AVDD.t1477 1.4705
R2242 AVDD.n1824 AVDD.t1448 1.4705
R2243 AVDD.n1819 AVDD.t1679 1.4705
R2244 AVDD.n1819 AVDD.t1589 1.4705
R2245 AVDD.n1814 AVDD.t1483 1.4705
R2246 AVDD.n1814 AVDD.t1645 1.4705
R2247 AVDD.n1812 AVDD.t1472 1.4705
R2248 AVDD.n1812 AVDD.t1454 1.4705
R2249 AVDD.n1913 AVDD.t1459 1.4705
R2250 AVDD.n1913 AVDD.t1465 1.4705
R2251 AVDD.n1914 AVDD.t1288 1.4705
R2252 AVDD.n1914 AVDD.t1295 1.4705
R2253 AVDD.n1907 AVDD.t1670 1.4705
R2254 AVDD.n1907 AVDD.t1684 1.4705
R2255 AVDD.n1908 AVDD.t1661 1.4705
R2256 AVDD.n1908 AVDD.t1675 1.4705
R2257 AVDD.n1649 AVDD.t1399 1.4705
R2258 AVDD.n1649 AVDD.t1581 1.4705
R2259 AVDD.n1657 AVDD.t1672 1.4705
R2260 AVDD.n1657 AVDD.t1492 1.4705
R2261 AVDD.n1715 AVDD.t1656 1.4705
R2262 AVDD.n1715 AVDD.t1590 1.4705
R2263 AVDD.n1716 AVDD.t1375 1.4705
R2264 AVDD.n1716 AVDD.t1649 1.4705
R2265 AVDD.n1718 AVDD.t1440 1.4705
R2266 AVDD.n1718 AVDD.t1387 1.4705
R2267 AVDD.n1719 AVDD.t1432 1.4705
R2268 AVDD.n1719 AVDD.t1489 1.4705
R2269 AVDD.n1722 AVDD.t1450 1.4705
R2270 AVDD.n1722 AVDD.t1569 1.4705
R2271 AVDD.n1723 AVDD.t1476 1.4705
R2272 AVDD.n1723 AVDD.t1690 1.4705
R2273 AVDD.n1726 AVDD.t1463 1.4705
R2274 AVDD.n1726 AVDD.t1680 1.4705
R2275 AVDD.n1727 AVDD.t1293 1.4705
R2276 AVDD.n1727 AVDD.t1592 1.4705
R2277 AVDD.n1731 AVDD.t1424 1.4705
R2278 AVDD.n1731 AVDD.t1397 1.4705
R2279 AVDD.n1732 AVDD.t1437 1.4705
R2280 AVDD.n1732 AVDD.t1383 1.4705
R2281 AVDD.n1735 AVDD.t1429 1.4705
R2282 AVDD.n1735 AVDD.t1485 1.4705
R2283 AVDD.n1736 AVDD.t1405 1.4705
R2284 AVDD.n1736 AVDD.t1451 1.4705
R2285 AVDD.n1739 AVDD.t1473 1.4705
R2286 AVDD.n1739 AVDD.t1468 1.4705
R2287 AVDD.n1740 AVDD.t1462 1.4705
R2288 AVDD.n1740 AVDD.t1303 1.4705
R2289 AVDD.n1743 AVDD.t1404 1.4705
R2290 AVDD.n1743 AVDD.t1563 1.4705
R2291 AVDD.n1744 AVDD.t1393 1.4705
R2292 AVDD.n1744 AVDD.t1682 1.4705
R2293 AVDD.n1682 AVDD.t1480 1.4705
R2294 AVDD.n1682 AVDD.t1490 1.4705
R2295 AVDD.n1683 AVDD.t1689 1.4705
R2296 AVDD.n1683 AVDD.t1428 1.4705
R2297 AVDD.n1685 AVDD.t1475 1.4705
R2298 AVDD.n1685 AVDD.t1660 1.4705
R2299 AVDD.n1686 AVDD.t1494 1.4705
R2300 AVDD.n1686 AVDD.t1479 1.4705
R2301 AVDD.n1689 AVDD.t1688 1.4705
R2302 AVDD.n1689 AVDD.t1410 1.4705
R2303 AVDD.n1690 AVDD.t1647 1.4705
R2304 AVDD.n1690 AVDD.t1658 1.4705
R2305 AVDD.n1693 AVDD.t1582 1.4705
R2306 AVDD.n1693 AVDD.t1391 1.4705
R2307 AVDD.n1694 AVDD.t1474 1.4705
R2308 AVDD.n1694 AVDD.t1406 1.4705
R2309 AVDD.n1678 AVDD.t1447 1.4705
R2310 AVDD.n1678 AVDD.t1664 1.4705
R2311 AVDD.n1679 AVDD.t1441 1.4705
R2312 AVDD.n1679 AVDD.t1466 1.4705
R2313 AVDD.n1674 AVDD.t1460 1.4705
R2314 AVDD.n1674 AVDD.t1566 1.4705
R2315 AVDD.n1675 AVDD.t1654 1.4705
R2316 AVDD.n1675 AVDD.t1641 1.4705
R2317 AVDD.n1670 AVDD.t1674 1.4705
R2318 AVDD.n1670 AVDD.t1593 1.4705
R2319 AVDD.n1671 AVDD.t1445 1.4705
R2320 AVDD.n1671 AVDD.t1438 1.4705
R2321 AVDD.n1666 AVDD.t1671 1.4705
R2322 AVDD.n1666 AVDD.t1403 1.4705
R2323 AVDD.n1667 AVDD.t1296 1.4705
R2324 AVDD.n1667 AVDD.t1469 1.4705
R2325 AVDD.n1752 AVDD.t1667 1.4705
R2326 AVDD.n1752 AVDD.t1289 1.4705
R2327 AVDD.n1749 AVDD.t1578 1.4705
R2328 AVDD.n1749 AVDD.t1586 1.4705
R2329 AVDD.n1643 AVDD.t1573 1.4705
R2330 AVDD.n1643 AVDD.t1413 1.4705
R2331 AVDD.n1639 AVDD.t1417 1.4705
R2332 AVDD.n1639 AVDD.t1458 1.4705
R2333 AVDD.n1702 AVDD.t1416 1.4705
R2334 AVDD.n1702 AVDD.t1425 1.4705
R2335 AVDD.n1699 AVDD.t1431 1.4705
R2336 AVDD.n1699 AVDD.t1488 1.4705
R2337 AVDD.t853 AVDD.n1964 1.4705
R2338 AVDD.n1964 AVDD.t1112 1.4705
R2339 AVDD.n1965 AVDD.t1242 1.4705
R2340 AVDD.n1965 AVDD.t853 1.4705
R2341 AVDD.t988 AVDD.n1969 1.4705
R2342 AVDD.n1969 AVDD.t1242 1.4705
R2343 AVDD.n1972 AVDD.t610 1.4705
R2344 AVDD.n1972 AVDD.t1024 1.4705
R2345 AVDD.t331 AVDD.n1300 1.4705
R2346 AVDD.n1300 AVDD.t610 1.4705
R2347 AVDD.t137 AVDD.n1305 1.4705
R2348 AVDD.n1305 AVDD.t154 1.4705
R2349 AVDD.n1306 AVDD.t549 1.4705
R2350 AVDD.n1306 AVDD.t137 1.4705
R2351 AVDD.t1056 AVDD.n1310 1.4705
R2352 AVDD.n1310 AVDD.t549 1.4705
R2353 AVDD.n31 AVDD.t189 1.4705
R2354 AVDD.t466 AVDD.n31 1.4705
R2355 AVDD.n29 AVDD.t618 1.4705
R2356 AVDD.t189 AVDD.n29 1.4705
R2357 AVDD.n28 AVDD.t341 1.4705
R2358 AVDD.t618 AVDD.n28 1.4705
R2359 AVDD.t1228 AVDD.n25 1.4705
R2360 AVDD.t376 AVDD.n25 1.4705
R2361 AVDD.t964 AVDD.n1298 1.4705
R2362 AVDD.n1298 AVDD.t1228 1.4705
R2363 AVDD.n1297 AVDD.t800 1.4705
R2364 AVDD.t813 AVDD.n1297 1.4705
R2365 AVDD.n1295 AVDD.t1174 1.4705
R2366 AVDD.t800 AVDD.n1295 1.4705
R2367 AVDD.n1294 AVDD.t412 1.4705
R2368 AVDD.t1174 AVDD.n1294 1.4705
R2369 AVDD.n500 AVDD.t1164 1.4705
R2370 AVDD.t736 AVDD.n500 1.4705
R2371 AVDD.n495 AVDD.t280 1.4705
R2372 AVDD.n495 AVDD.t1164 1.4705
R2373 AVDD.n494 AVDD.t699 1.4705
R2374 AVDD.t280 AVDD.n494 1.4705
R2375 AVDD.n489 AVDD.t1234 1.4705
R2376 AVDD.t970 AVDD.n489 1.4705
R2377 AVDD.n484 AVDD.t382 1.4705
R2378 AVDD.n484 AVDD.t1234 1.4705
R2379 AVDD.n481 AVDD.t624 1.4705
R2380 AVDD.t348 AVDD.n481 1.4705
R2381 AVDD.n476 AVDD.t940 1.4705
R2382 AVDD.n476 AVDD.t624 1.4705
R2383 AVDD.n475 AVDD.t1200 1.4705
R2384 AVDD.t940 AVDD.n475 1.4705
R2385 AVDD.n498 AVDD.t292 1.4705
R2386 AVDD.n498 AVDD.t1140 1.4705
R2387 AVDD.n497 AVDD.t675 1.4705
R2388 AVDD.t292 AVDD.n497 1.4705
R2389 AVDD.n492 AVDD.t1078 1.4705
R2390 AVDD.n492 AVDD.t675 1.4705
R2391 AVDD.n487 AVDD.t364 1.4705
R2392 AVDD.n487 AVDD.t60 1.4705
R2393 AVDD.n486 AVDD.t804 1.4705
R2394 AVDD.t364 AVDD.n486 1.4705
R2395 AVDD.n479 AVDD.t1022 1.4705
R2396 AVDD.n479 AVDD.t758 1.4705
R2397 AVDD.n478 AVDD.t20 1.4705
R2398 AVDD.t1022 AVDD.n478 1.4705
R2399 AVDD.n473 AVDD.t333 1.4705
R2400 AVDD.n473 AVDD.t20 1.4705
R2401 AVDD.t120 AVDD.n413 1.4705
R2402 AVDD.n413 AVDD.t558 1.4705
R2403 AVDD.n414 AVDD.t400 1.4705
R2404 AVDD.n414 AVDD.t120 1.4705
R2405 AVDD.t839 AVDD.n418 1.4705
R2406 AVDD.n418 AVDD.t400 1.4705
R2407 AVDD.n421 AVDD.t1052 1.4705
R2408 AVDD.n421 AVDD.t796 1.4705
R2409 AVDD.t201 AVDD.n426 1.4705
R2410 AVDD.n426 AVDD.t1052 1.4705
R2411 AVDD.t505 AVDD.n431 1.4705
R2412 AVDD.n431 AVDD.t227 1.4705
R2413 AVDD.n432 AVDD.t1030 1.4705
R2414 AVDD.n432 AVDD.t505 1.4705
R2415 AVDD.t1280 AVDD.n436 1.4705
R2416 AVDD.n436 AVDD.t1030 1.4705
R2417 AVDD.n410 AVDD.t523 1.4705
R2418 AVDD.n410 AVDD.t950 1.4705
R2419 AVDD.n408 AVDD.t815 1.4705
R2420 AVDD.t523 AVDD.n408 1.4705
R2421 AVDD.n407 AVDD.t1218 1.4705
R2422 AVDD.t815 AVDD.n407 1.4705
R2423 AVDD.n404 AVDD.t176 1.4705
R2424 AVDD.t1176 AVDD.n404 1.4705
R2425 AVDD.n403 AVDD.t612 1.4705
R2426 AVDD.t176 AVDD.n403 1.4705
R2427 AVDD.n401 AVDD.t916 1.4705
R2428 AVDD.t630 AVDD.n401 1.4705
R2429 AVDD.n399 AVDD.t149 1.4705
R2430 AVDD.t916 AVDD.n399 1.4705
R2431 AVDD.n398 AVDD.t434 1.4705
R2432 AVDD.t149 AVDD.n398 1.4705
R2433 AVDD.t1040 AVDD.n1381 1.4705
R2434 AVDD.n1381 AVDD.t454 1.4705
R2435 AVDD.n1382 AVDD.t1110 1.4705
R2436 AVDD.n1382 AVDD.t1040 1.4705
R2437 AVDD.t762 AVDD.n1386 1.4705
R2438 AVDD.n1386 AVDD.t1110 1.4705
R2439 AVDD.n1389 AVDD.t231 1.4705
R2440 AVDD.n1389 AVDD.t157 1.4705
R2441 AVDD.n614 AVDD.t1146 1.4705
R2442 AVDD.t231 AVDD.n614 1.4705
R2443 AVDD.n609 AVDD.t535 1.4705
R2444 AVDD.t462 AVDD.n609 1.4705
R2445 AVDD.n604 AVDD.t165 1.4705
R2446 AVDD.n604 AVDD.t535 1.4705
R2447 AVDD.n603 AVDD.t244 1.4705
R2448 AVDD.t165 AVDD.n603 1.4705
R2449 AVDD.n593 AVDD.t786 1.4705
R2450 AVDD.t1148 AVDD.n593 1.4705
R2451 AVDD.n588 AVDD.t857 1.4705
R2452 AVDD.n588 AVDD.t786 1.4705
R2453 AVDD.n587 AVDD.t460 1.4705
R2454 AVDD.t857 AVDD.n587 1.4705
R2455 AVDD.n582 AVDD.t908 1.4705
R2456 AVDD.t859 AVDD.n582 1.4705
R2457 AVDD.n577 AVDD.t531 1.4705
R2458 AVDD.n577 AVDD.t908 1.4705
R2459 AVDD.n574 AVDD.t1270 1.4705
R2460 AVDD.t1224 AVDD.n574 1.4705
R2461 AVDD.n569 AVDD.t768 1.4705
R2462 AVDD.n569 AVDD.t1270 1.4705
R2463 AVDD.n568 AVDD.t821 1.4705
R2464 AVDD.t768 AVDD.n568 1.4705
R2465 AVDD.n619 AVDD.t1048 1.4705
R2466 AVDD.t464 AVDD.n619 1.4705
R2467 AVDD.n617 AVDD.t1118 1.4705
R2468 AVDD.t1048 AVDD.n617 1.4705
R2469 AVDD.n616 AVDD.t770 1.4705
R2470 AVDD.t1118 AVDD.n616 1.4705
R2471 AVDD.t236 AVDD.n115 1.4705
R2472 AVDD.t161 AVDD.n115 1.4705
R2473 AVDD.t1152 AVDD.n611 1.4705
R2474 AVDD.n611 AVDD.t236 1.4705
R2475 AVDD.n607 AVDD.t541 1.4705
R2476 AVDD.n607 AVDD.t474 1.4705
R2477 AVDD.n606 AVDD.t173 1.4705
R2478 AVDD.t541 AVDD.n606 1.4705
R2479 AVDD.n601 AVDD.t250 1.4705
R2480 AVDD.n601 AVDD.t173 1.4705
R2481 AVDD.n591 AVDD.t788 1.4705
R2482 AVDD.n591 AVDD.t1156 1.4705
R2483 AVDD.n590 AVDD.t865 1.4705
R2484 AVDD.t788 AVDD.n590 1.4705
R2485 AVDD.n585 AVDD.t468 1.4705
R2486 AVDD.n585 AVDD.t865 1.4705
R2487 AVDD.n580 AVDD.t914 1.4705
R2488 AVDD.n580 AVDD.t861 1.4705
R2489 AVDD.n579 AVDD.t539 1.4705
R2490 AVDD.t914 AVDD.n579 1.4705
R2491 AVDD.n572 AVDD.t1274 1.4705
R2492 AVDD.n572 AVDD.t1230 1.4705
R2493 AVDD.n571 AVDD.t772 1.4705
R2494 AVDD.t1274 AVDD.n571 1.4705
R2495 AVDD.n566 AVDD.t829 1.4705
R2496 AVDD.n566 AVDD.t772 1.4705
R2497 AVDD.t689 AVDD.n521 1.4705
R2498 AVDD.n521 AVDD.t275 1.4705
R2499 AVDD.n522 AVDD.t1062 1.4705
R2500 AVDD.n522 AVDD.t689 1.4705
R2501 AVDD.t218 AVDD.n526 1.4705
R2502 AVDD.n526 AVDD.t1062 1.4705
R2503 AVDD.n529 AVDD.t792 1.4705
R2504 AVDD.n529 AVDD.t491 1.4705
R2505 AVDD.t1190 AVDD.n534 1.4705
R2506 AVDD.n534 AVDD.t792 1.4705
R2507 AVDD.t134 AVDD.n539 1.4705
R2508 AVDD.n539 AVDD.t1160 1.4705
R2509 AVDD.n540 AVDD.t446 1.4705
R2510 AVDD.n540 AVDD.t134 1.4705
R2511 AVDD.t750 AVDD.n544 1.4705
R2512 AVDD.n544 AVDD.t446 1.4705
R2513 AVDD.t944 AVDD.n372 1.4705
R2514 AVDD.n372 AVDD.t51 1.4705
R2515 AVDD.n373 AVDD.t1202 1.4705
R2516 AVDD.n373 AVDD.t944 1.4705
R2517 AVDD.t360 AVDD.n377 1.4705
R2518 AVDD.n377 AVDD.t1202 1.4705
R2519 AVDD.n380 AVDD.t590 1.4705
R2520 AVDD.n380 AVDD.t317 1.4705
R2521 AVDD.t1012 AVDD.n385 1.4705
R2522 AVDD.n385 AVDD.t590 1.4705
R2523 AVDD.t1278 AVDD.n390 1.4705
R2524 AVDD.n390 AVDD.t1028 1.4705
R2525 AVDD.n391 AVDD.t580 1.4705
R2526 AVDD.n391 AVDD.t1278 1.4705
R2527 AVDD.t873 AVDD.n395 1.4705
R2528 AVDD.n395 AVDD.t580 1.4705
R2529 AVDD.t661 AVDD.n1422 1.4705
R2530 AVDD.n1422 AVDD.t242 1.4705
R2531 AVDD.n1423 AVDD.t1034 1.4705
R2532 AVDD.n1423 AVDD.t661 1.4705
R2533 AVDD.t194 AVDD.n1427 1.4705
R2534 AVDD.n1427 AVDD.t1034 1.4705
R2535 AVDD.n1430 AVDD.t764 1.4705
R2536 AVDD.n1430 AVDD.t456 1.4705
R2537 AVDD.t1172 AVDD.n330 1.4705
R2538 AVDD.n330 AVDD.t764 1.4705
R2539 AVDD.t123 AVDD.n335 1.4705
R2540 AVDD.n335 AVDD.t1128 1.4705
R2541 AVDD.n336 AVDD.t424 1.4705
R2542 AVDD.n336 AVDD.t123 1.4705
R2543 AVDD.t728 AVDD.n340 1.4705
R2544 AVDD.n340 AVDD.t424 1.4705
R2545 AVDD.n100 AVDD.t1268 1.4705
R2546 AVDD.t886 AVDD.n100 1.4705
R2547 AVDD.n98 AVDD.t404 1.4705
R2548 AVDD.t1268 AVDD.n98 1.4705
R2549 AVDD.n97 AVDD.t847 1.4705
R2550 AVDD.t404 AVDD.n97 1.4705
R2551 AVDD.t89 AVDD.n94 1.4705
R2552 AVDD.t1092 AVDD.n94 1.4705
R2553 AVDD.t525 AVDD.n328 1.4705
R2554 AVDD.n328 AVDD.t89 1.4705
R2555 AVDD.n327 AVDD.t778 1.4705
R2556 AVDD.t483 AVDD.n327 1.4705
R2557 AVDD.n325 AVDD.t1058 1.4705
R2558 AVDD.t778 AVDD.n325 1.4705
R2559 AVDD.n324 AVDD.t45 1.4705
R2560 AVDD.t1058 AVDD.n324 1.4705
R2561 AVDD.n1450 AVDD.t780 1.4705
R2562 AVDD.t345 AVDD.n1450 1.4705
R2563 AVDD.n1446 AVDD.t1162 1.4705
R2564 AVDD.n1446 AVDD.t780 1.4705
R2565 AVDD.n1445 AVDD.t307 1.4705
R2566 AVDD.t1162 AVDD.n1445 1.4705
R2567 AVDD.n1440 AVDD.t871 1.4705
R2568 AVDD.t576 AVDD.n1440 1.4705
R2569 AVDD.t1254 AVDD.n298 1.4705
R2570 AVDD.n298 AVDD.t871 1.4705
R2571 AVDD.t224 AVDD.n303 1.4705
R2572 AVDD.n303 AVDD.t1214 1.4705
R2573 AVDD.n304 AVDD.t537 1.4705
R2574 AVDD.n304 AVDD.t224 1.4705
R2575 AVDD.t827 AVDD.n308 1.4705
R2576 AVDD.n308 AVDD.t537 1.4705
R2577 AVDD.n1537 AVDD.t1308 1.4705
R2578 AVDD.n1537 AVDD.t1634 1.4705
R2579 AVDD.n1538 AVDD.t1317 1.4705
R2580 AVDD.n1538 AVDD.t1560 1.4705
R2581 AVDD.n1487 AVDD.t1354 1.4705
R2582 AVDD.n1487 AVDD.t1608 1.4705
R2583 AVDD.n1488 AVDD.t1522 1.4705
R2584 AVDD.n1488 AVDD.t1615 1.4705
R2585 AVDD.n1597 AVDD.t1502 1.4705
R2586 AVDD.n1597 AVDD.t1320 1.4705
R2587 AVDD.n1595 AVDD.t1350 1.4705
R2588 AVDD.n1595 AVDD.t1338 1.4705
R2589 AVDD.n1593 AVDD.t1325 1.4705
R2590 AVDD.n1593 AVDD.t1629 1.4705
R2591 AVDD.n1591 AVDD.t1513 1.4705
R2592 AVDD.n1591 AVDD.t1547 1.4705
R2593 AVDD.n75 AVDD.t1531 1.4705
R2594 AVDD.n75 AVDD.t1365 1.4705
R2595 AVDD.n73 AVDD.t1370 1.4705
R2596 AVDD.n73 AVDD.t1625 1.4705
R2597 AVDD.n71 AVDD.t1309 1.4705
R2598 AVDD.n71 AVDD.t1614 1.4705
R2599 AVDD.n70 AVDD.t1527 1.4705
R2600 AVDD.n70 AVDD.t1339 1.4705
R2601 AVDD.n1484 AVDD.t1621 1.4705
R2602 AVDD.n1484 AVDD.t1368 1.4705
R2603 AVDD.n1481 AVDD.t1553 1.4705
R2604 AVDD.n1481 AVDD.t1315 1.4705
R2605 AVDD.n1478 AVDD.t1372 1.4705
R2606 AVDD.n1478 AVDD.t1606 1.4705
R2607 AVDD.n1475 AVDD.t1632 1.4705
R2608 AVDD.n1475 AVDD.t1376 1.4705
R2609 AVDD.n1470 AVDD.t1514 1.4705
R2610 AVDD.n1470 AVDD.t1343 1.4705
R2611 AVDD.n1465 AVDD.t1347 1.4705
R2612 AVDD.n1465 AVDD.t1336 1.4705
R2613 AVDD.n1460 AVDD.t1357 1.4705
R2614 AVDD.n1460 AVDD.t1326 1.4705
R2615 AVDD.n1458 AVDD.t1506 1.4705
R2616 AVDD.n1458 AVDD.t1541 1.4705
R2617 AVDD.n1558 AVDD.t1305 1.4705
R2618 AVDD.n1558 AVDD.t1542 1.4705
R2619 AVDD.n1556 AVDD.t1509 1.4705
R2620 AVDD.n1556 AVDD.t1559 1.4705
R2621 AVDD.n1554 AVDD.t1550 1.4705
R2622 AVDD.n1554 AVDD.t1362 1.4705
R2623 AVDD.n1552 AVDD.t1314 1.4705
R2624 AVDD.n1552 AVDD.t1618 1.4705
R2625 AVDD.n1549 AVDD.t1337 1.4705
R2626 AVDD.n1549 AVDD.t1518 1.4705
R2627 AVDD.n1547 AVDD.t1523 1.4705
R2628 AVDD.n1547 AVDD.t1355 1.4705
R2629 AVDD.n1545 AVDD.t1532 1.4705
R2630 AVDD.n1545 AVDD.t1345 1.4705
R2631 AVDD.n1544 AVDD.t1331 1.4705
R2632 AVDD.n1544 AVDD.t1638 1.4705
R2633 AVDD.n1521 AVDD.t1610 1.4705
R2634 AVDD.n1521 AVDD.t1546 1.4705
R2635 AVDD.n1518 AVDD.t1512 1.4705
R2636 AVDD.n1518 AVDD.t1335 1.4705
R2637 AVDD.n1515 AVDD.t1535 1.4705
R2638 AVDD.n1515 AVDD.t1543 1.4705
R2639 AVDD.n1512 AVDD.t1349 1.4705
R2640 AVDD.n1512 AVDD.t1359 1.4705
R2641 AVDD.n1507 AVDD.t1508 1.4705
R2642 AVDD.n1507 AVDD.t1332 1.4705
R2643 AVDD.n1502 AVDD.t1544 1.4705
R2644 AVDD.n1502 AVDD.t1498 1.4705
R2645 AVDD.n1497 AVDD.t1311 1.4705
R2646 AVDD.n1497 AVDD.t1319 1.4705
R2647 AVDD.n1495 AVDD.t1501 1.4705
R2648 AVDD.n1495 AVDD.t1511 1.4705
R2649 AVDD.n1583 AVDD.t1505 1.4705
R2650 AVDD.n1583 AVDD.t1556 1.4705
R2651 AVDD.n1584 AVDD.t1495 1.4705
R2652 AVDD.n1584 AVDD.t1551 1.4705
R2653 AVDD.n1576 AVDD.t1622 1.4705
R2654 AVDD.n1576 AVDD.t1534 1.4705
R2655 AVDD.n1577 AVDD.t1612 1.4705
R2656 AVDD.n1577 AVDD.t1526 1.4705
R2657 AVDD.n207 AVDD.t1352 1.4705
R2658 AVDD.n207 AVDD.t1361 1.4705
R2659 AVDD.n201 AVDD.t1630 1.4705
R2660 AVDD.n201 AVDD.t1497 1.4705
R2661 AVDD.n272 AVDD.t1516 1.4705
R2662 AVDD.n272 AVDD.t1334 1.4705
R2663 AVDD.n273 AVDD.t1507 1.4705
R2664 AVDD.n273 AVDD.t1323 1.4705
R2665 AVDD.n275 AVDD.t1367 1.4705
R2666 AVDD.n275 AVDD.t1620 1.4705
R2667 AVDD.n276 AVDD.t1356 1.4705
R2668 AVDD.n276 AVDD.t1609 1.4705
R2669 AVDD.n279 AVDD.t1605 1.4705
R2670 AVDD.n279 AVDD.t1503 1.4705
R2671 AVDD.n280 AVDD.t1329 1.4705
R2672 AVDD.n280 AVDD.t1635 1.4705
R2673 AVDD.n283 AVDD.t1525 1.4705
R2674 AVDD.n283 AVDD.t1561 1.4705
R2675 AVDD.n284 AVDD.t1517 1.4705
R2676 AVDD.n284 AVDD.t1552 1.4705
R2677 AVDD.n268 AVDD.t1548 1.4705
R2678 AVDD.n268 AVDD.t1310 1.4705
R2679 AVDD.n269 AVDD.t1538 1.4705
R2680 AVDD.n269 AVDD.t1369 1.4705
R2681 AVDD.n264 AVDD.t1313 1.4705
R2682 AVDD.n264 AVDD.t1499 1.4705
R2683 AVDD.n265 AVDD.t1306 1.4705
R2684 AVDD.n265 AVDD.t1627 1.4705
R2685 AVDD.n260 AVDD.t1324 1.4705
R2686 AVDD.n260 AVDD.t1628 1.4705
R2687 AVDD.n261 AVDD.t1312 1.4705
R2688 AVDD.n261 AVDD.t1617 1.4705
R2689 AVDD.n256 AVDD.t1540 1.4705
R2690 AVDD.n256 AVDD.t1353 1.4705
R2691 AVDD.n257 AVDD.t1528 1.4705
R2692 AVDD.n257 AVDD.t1342 1.4705
R2693 AVDD.n180 AVDD.t1321 1.4705
R2694 AVDD.n180 AVDD.t1554 1.4705
R2695 AVDD.n181 AVDD.t1328 1.4705
R2696 AVDD.n181 AVDD.t1530 1.4705
R2697 AVDD.n183 AVDD.t1519 1.4705
R2698 AVDD.n183 AVDD.t1351 1.4705
R2699 AVDD.n184 AVDD.t1496 1.4705
R2700 AVDD.n184 AVDD.t1322 1.4705
R2701 AVDD.n187 AVDD.t1340 1.4705
R2702 AVDD.n187 AVDD.t1307 1.4705
R2703 AVDD.n188 AVDD.t1521 1.4705
R2704 AVDD.n188 AVDD.t1378 1.4705
R2705 AVDD.n191 AVDD.t1330 1.4705
R2706 AVDD.n191 AVDD.t1637 1.4705
R2707 AVDD.n192 AVDD.t1558 1.4705
R2708 AVDD.n192 AVDD.t1344 1.4705
R2709 AVDD.n214 AVDD.t1619 1.4705
R2710 AVDD.n214 AVDD.t1533 1.4705
R2711 AVDD.n215 AVDD.t1636 1.4705
R2712 AVDD.n215 AVDD.t1316 1.4705
R2713 AVDD.n218 AVDD.t1539 1.4705
R2714 AVDD.n218 AVDD.t1371 1.4705
R2715 AVDD.n219 AVDD.t1529 1.4705
R2716 AVDD.n219 AVDD.t1624 1.4705
R2717 AVDD.n222 AVDD.t1549 1.4705
R2718 AVDD.n222 AVDD.t1360 1.4705
R2719 AVDD.n223 AVDD.t1366 1.4705
R2720 AVDD.n223 AVDD.t1304 1.4705
R2721 AVDD.n226 AVDD.t1613 1.4705
R2722 AVDD.n226 AVDD.t1510 1.4705
R2723 AVDD.n227 AVDD.t1626 1.4705
R2724 AVDD.n227 AVDD.t1639 1.4705
R2725 AVDD.n144 AVDD.t1633 1.4705
R2726 AVDD.n144 AVDD.t1545 1.4705
R2727 AVDD.n292 AVDD.t1607 1.4705
R2728 AVDD.n292 AVDD.t1520 1.4705
R2729 AVDD.n250 AVDD.t1524 1.4705
R2730 AVDD.n250 AVDD.t1557 1.4705
R2731 AVDD.n244 AVDD.t1500 1.4705
R2732 AVDD.n244 AVDD.t1536 1.4705
R2733 AVDD.n231 AVDD.t1364 1.4705
R2734 AVDD.n231 AVDD.t1616 1.4705
R2735 AVDD.n235 AVDD.t1341 1.4705
R2736 AVDD.n235 AVDD.t1327 1.4705
R2737 AVDD.n1350 AVDD.t918 1.4705
R2738 AVDD.t23 AVDD.n1350 1.4705
R2739 AVDD.n1345 AVDD.t1182 1.4705
R2740 AVDD.n1345 AVDD.t918 1.4705
R2741 AVDD.n1344 AVDD.t339 1.4705
R2742 AVDD.t1182 AVDD.n1344 1.4705
R2743 AVDD.n1339 AVDD.t568 1.4705
R2744 AVDD.t299 AVDD.n1339 1.4705
R2745 AVDD.n1334 AVDD.t994 1.4705
R2746 AVDD.n1334 AVDD.t568 1.4705
R2747 AVDD.n1331 AVDD.t1266 1.4705
R2748 AVDD.t1010 AVDD.n1331 1.4705
R2749 AVDD.n1326 AVDD.t560 1.4705
R2750 AVDD.n1326 AVDD.t1266 1.4705
R2751 AVDD.n1325 AVDD.t845 1.4705
R2752 AVDD.t560 AVDD.n1325 1.4705
R2753 AVDD.n1348 AVDD.t277 1.4705
R2754 AVDD.n1348 AVDD.t693 1.4705
R2755 AVDD.n1347 AVDD.t553 1.4705
R2756 AVDD.t277 AVDD.n1347 1.4705
R2757 AVDD.n1342 AVDD.t974 1.4705
R2758 AVDD.n1342 AVDD.t553 1.4705
R2759 AVDD.n1337 AVDD.t1194 1.4705
R2760 AVDD.n1337 AVDD.t928 1.4705
R2761 AVDD.n1336 AVDD.t352 1.4705
R2762 AVDD.t1194 AVDD.n1336 1.4705
R2763 AVDD.n1329 AVDD.t649 1.4705
R2764 AVDD.n1329 AVDD.t369 1.4705
R2765 AVDD.n1328 AVDD.t1180 1.4705
R2766 AVDD.t649 AVDD.n1328 1.4705
R2767 AVDD.n1323 AVDD.t179 1.4705
R2768 AVDD.n1323 AVDD.t1180 1.4705
R2769 AVDD.n1141 AVDD.t1186 1.4705
R2770 AVDD.n1141 AVDD.t790 1.4705
R2771 AVDD.n1140 AVDD.t922 1.4705
R2772 AVDD.t1186 AVDD.n1140 1.4705
R2773 AVDD.t216 AVDD.n718 1.4705
R2774 AVDD.n718 AVDD.t641 1.4705
R2775 AVDD.n719 AVDD.t273 1.4705
R2776 AVDD.n719 AVDD.t216 1.4705
R2777 AVDD.t65 AVDD.n891 1.4705
R2778 AVDD.n891 AVDD.t511 1.4705
R2779 AVDD.n892 AVDD.t657 1.4705
R2780 AVDD.n892 AVDD.t65 1.4705
R2781 AVDD.n882 AVDD.t229 1.4705
R2782 AVDD.n882 AVDD.t657 1.4705
R2783 AVDD.n865 AVDD.t880 1.4705
R2784 AVDD.t1154 AVDD.n865 1.4705
R2785 AVDD.n713 AVDD.t744 1.4705
R2786 AVDD.n713 AVDD.t1204 1.4705
R2787 AVDD.n708 AVDD.t367 1.4705
R2788 AVDD.t744 AVDD.n708 1.4705
R2789 AVDD.t1252 AVDD.n722 1.4705
R2790 AVDD.n722 AVDD.t367 1.4705
R2791 AVDD.n886 AVDD.t1122 1.4705
R2792 AVDD.t1044 AVDD.n886 1.4705
R2793 AVDD.n885 AVDD.t28 1.4705
R2794 AVDD.t1122 AVDD.n885 1.4705
R2795 AVDD.n879 AVDD.t902 1.4705
R2796 AVDD.t687 AVDD.n879 1.4705
R2797 AVDD.n873 AVDD.t962 1.4705
R2798 AVDD.n873 AVDD.t902 1.4705
R2799 AVDD.n872 AVDD.t476 1.4705
R2800 AVDD.t962 AVDD.n872 1.4705
R2801 AVDD.n1145 AVDD.t790 1.4705
R2802 AVDD.t740 AVDD.n1145 1.4705
R2803 AVDD.n861 AVDD.t1260 1.4705
R2804 AVDD.t880 AVDD.n861 1.4705
R2805 AVDD.n855 AVDD.t1006 1.4705
R2806 AVDD.n855 AVDD.t1260 1.4705
R2807 AVDD.n852 AVDD.t632 1.4705
R2808 AVDD.t1042 AVDD.n852 1.4705
R2809 AVDD.t356 AVDD.n1981 1.4705
R2810 AVDD.n1981 AVDD.t632 1.4705
R2811 AVDD.t171 AVDD.n1986 1.4705
R2812 AVDD.n1986 AVDD.t184 1.4705
R2813 AVDD.n1987 AVDD.t572 1.4705
R2814 AVDD.n1987 AVDD.t171 1.4705
R2815 AVDD.t1074 AVDD.n1991 1.4705
R2816 AVDD.n1991 AVDD.t572 1.4705
R2817 AVDD.n820 AVDD.t31 1.4705
R2818 AVDD.t336 AVDD.n820 1.4705
R2819 AVDD.n815 AVDD.t470 1.4705
R2820 AVDD.n815 AVDD.t31 1.4705
R2821 AVDD.n814 AVDD.t196 1.4705
R2822 AVDD.t470 AVDD.n814 1.4705
R2823 AVDD.n809 AVDD.t1086 1.4705
R2824 AVDD.t253 AVDD.n809 1.4705
R2825 AVDD.n804 AVDD.t835 1.4705
R2826 AVDD.n804 AVDD.t1086 1.4705
R2827 AVDD.n801 AVDD.t645 1.4705
R2828 AVDD.t663 AVDD.n801 1.4705
R2829 AVDD.n796 AVDD.t1026 1.4705
R2830 AVDD.n796 AVDD.t645 1.4705
R2831 AVDD.n795 AVDD.t295 1.4705
R2832 AVDD.t1026 AVDD.n795 1.4705
R2833 AVDD.n818 AVDD.t444 1.4705
R2834 AVDD.n818 AVDD.t746 1.4705
R2835 AVDD.n817 AVDD.t892 1.4705
R2836 AVDD.t444 AVDD.n817 1.4705
R2837 AVDD.n812 AVDD.t602 1.4705
R2838 AVDD.n812 AVDD.t892 1.4705
R2839 AVDD.n807 AVDD.t220 1.4705
R2840 AVDD.n807 AVDD.t647 1.4705
R2841 AVDD.n806 AVDD.t1212 1.4705
R2842 AVDD.t220 AVDD.n806 1.4705
R2843 AVDD.n799 AVDD.t1032 1.4705
R2844 AVDD.n799 AVDD.t1054 1.4705
R2845 AVDD.n798 AVDD.t142 1.4705
R2846 AVDD.t1032 AVDD.n798 1.4705
R2847 AVDD.n793 AVDD.t683 1.4705
R2848 AVDD.n793 AVDD.t142 1.4705
R2849 AVDD.t1232 AVDD.n756 1.4705
R2850 AVDD.n756 AVDD.t1198 1.4705
R2851 AVDD.n757 AVDD.t379 1.4705
R2852 AVDD.n757 AVDD.t1232 1.4705
R2853 AVDD.t94 AVDD.n761 1.4705
R2854 AVDD.n761 AVDD.t379 1.4705
R2855 AVDD.n764 AVDD.t697 1.4705
R2856 AVDD.n764 AVDD.t1102 1.4705
R2857 AVDD.t734 AVDD.n769 1.4705
R2858 AVDD.n769 AVDD.t697 1.4705
R2859 AVDD.t562 AVDD.n774 1.4705
R2860 AVDD.n774 AVDD.t986 1.4705
R2861 AVDD.n775 AVDD.t1124 1.4705
R2862 AVDD.n775 AVDD.t562 1.4705
R2863 AVDD.t709 AVDD.n779 1.4705
R2864 AVDD.n779 AVDD.t1124 1.4705
R2865 AVDD.n742 AVDD.t362 1.4705
R2866 AVDD.t326 AVDD.n742 1.4705
R2867 AVDD.n740 AVDD.t802 1.4705
R2868 AVDD.t362 AVDD.n740 1.4705
R2869 AVDD.n739 AVDD.t507 1.4705
R2870 AVDD.t802 AVDD.n739 1.4705
R2871 AVDD.n736 AVDD.t1072 1.4705
R2872 AVDD.t234 AVDD.n736 1.4705
R2873 AVDD.n735 AVDD.t1138 1.4705
R2874 AVDD.t1072 AVDD.n735 1.4705
R2875 AVDD.n733 AVDD.t956 1.4705
R2876 AVDD.t83 AVDD.n733 1.4705
R2877 AVDD.n731 AVDD.t256 1.4705
R2878 AVDD.t956 AVDD.n731 1.4705
R2879 AVDD.n730 AVDD.t1088 1.4705
R2880 AVDD.t256 AVDD.n730 1.4705
R2881 AVDD.n1133 AVDD.t1599 1.4705
R2882 AVDD.n1133 AVDD.t1285 1.4705
R2883 AVDD.n1131 AVDD.t1691 1.4705
R2884 AVDD.n1131 AVDD.t1696 1.4705
R2885 AVDD.n1128 AVDD.t1390 1.4705
R2886 AVDD.n1128 AVDD.t1434 1.4705
R2887 AVDD.n1126 AVDD.t1603 1.4705
R2888 AVDD.n1126 AVDD.t1597 1.4705
R2889 AVDD.n1124 AVDD.t1697 1.4705
R2890 AVDD.n1124 AVDD.t1604 1.4705
R2891 AVDD.n681 AVDD.t1407 1.4705
R2892 AVDD.n681 AVDD.t1298 1.4705
R2893 AVDD.n678 AVDD.t1287 1.4705
R2894 AVDD.n678 AVDD.t1595 1.4705
R2895 AVDD.n675 AVDD.t1471 1.4705
R2896 AVDD.n675 AVDD.t1444 1.4705
R2897 AVDD.n670 AVDD.t1380 1.4705
R2898 AVDD.n670 AVDD.t1412 1.4705
R2899 AVDD.n667 AVDD.t1646 1.4705
R2900 AVDD.n667 AVDD.t1481 1.4705
R2901 AVDD.n1091 AVDD.t1290 1.4705
R2902 AVDD.n1091 AVDD.t1651 1.4705
R2903 AVDD.n1093 AVDD.t1585 1.4705
R2904 AVDD.n1093 AVDD.t1382 1.4705
R2905 AVDD.n1085 AVDD.t1426 1.4705
R2906 AVDD.n1085 AVDD.t1381 1.4705
R2907 AVDD.n1087 AVDD.t1486 1.4705
R2908 AVDD.n1087 AVDD.t1666 1.4705
R2909 AVDD.n1079 AVDD.t1602 1.4705
R2910 AVDD.n1079 AVDD.t1600 1.4705
R2911 AVDD.n1081 AVDD.t1692 1.4705
R2912 AVDD.n1081 AVDD.t1284 1.4705
R2913 AVDD.n1069 AVDD.t1575 1.4705
R2914 AVDD.n1069 AVDD.t1302 1.4705
R2915 AVDD.n1071 AVDD.t1418 1.4705
R2916 AVDD.n1071 AVDD.t1677 1.4705
R2917 AVDD.n1063 AVDD.t1455 1.4705
R2918 AVDD.n1063 AVDD.t1565 1.4705
R2919 AVDD.n1065 AVDD.t1574 1.4705
R2920 AVDD.n1065 AVDD.t1436 1.4705
R2921 AVDD.n947 AVDD.t1291 1.4705
R2922 AVDD.n947 AVDD.t1653 1.4705
R2923 AVDD.n949 AVDD.t1640 1.4705
R2924 AVDD.n949 AVDD.t1384 1.4705
R2925 AVDD.n952 AVDD.t1415 1.4705
R2926 AVDD.n952 AVDD.t1676 1.4705
R2927 AVDD.n954 AVDD.t1576 1.4705
R2928 AVDD.n954 AVDD.t1461 1.4705
R2929 AVDD.n956 AVDD.t1457 1.4705
R2930 AVDD.n956 AVDD.t1568 1.4705
R2931 AVDD.n916 AVDD.t1699 1.4705
R2932 AVDD.n916 AVDD.t1281 1.4705
R2933 AVDD.n913 AVDD.t1283 1.4705
R2934 AVDD.n913 AVDD.t1693 1.4705
R2935 AVDD.n910 AVDD.t1650 1.4705
R2936 AVDD.n910 AVDD.t1587 1.4705
R2937 AVDD.n905 AVDD.t1598 1.4705
R2938 AVDD.n905 AVDD.t1698 1.4705
R2939 AVDD.n902 AVDD.t1695 1.4705
R2940 AVDD.n902 AVDD.t1601 1.4705
R2941 AVDD.n1024 AVDD.t324 1.4705
R2942 AVDD.t811 AVDD.n1024 1.4705
R2943 AVDD.n1020 AVDD.t1222 1.4705
R2944 AVDD.n1020 AVDD.t324 1.4705
R2945 AVDD.n1019 AVDD.t876 1.4705
R2946 AVDD.t1222 AVDD.n1019 1.4705
R2947 AVDD.n1014 AVDD.t718 1.4705
R2948 AVDD.t639 AVDD.n1014 1.4705
R2949 AVDD.n1009 AVDD.t926 1.4705
R2950 AVDD.n1009 AVDD.t718 1.4705
R2951 AVDD.n1006 AVDD.t481 1.4705
R2952 AVDD.t283 AVDD.n1006 1.4705
R2953 AVDD.n1002 AVDD.t556 1.4705
R2954 AVDD.n1002 AVDD.t481 1.4705
R2955 AVDD.n1001 AVDD.t40 1.4705
R2956 AVDD.t556 AVDD.n1001 1.4705
R2957 AVDD.n1198 AVDD.t86 1.4705
R2958 AVDD.n1198 AVDD.t34 1.4705
R2959 AVDD.n1197 AVDD.t519 1.4705
R2960 AVDD.t86 AVDD.n1197 1.4705
R2961 AVDD.n1192 AVDD.t258 1.4705
R2962 AVDD.n1192 AVDD.t519 1.4705
R2963 AVDD.n1187 AVDD.t841 1.4705
R2964 AVDD.n1187 AVDD.t1240 1.4705
R2965 AVDD.n1186 AVDD.t884 1.4705
R2966 AVDD.t841 AVDD.n1186 1.4705
R2967 AVDD.n1179 AVDD.t705 1.4705
R2968 AVDD.n1179 AVDD.t1114 1.4705
R2969 AVDD.n1178 AVDD.t1244 1.4705
R2970 AVDD.t705 AVDD.n1178 1.4705
R2971 AVDD.n1173 AVDD.t851 1.4705
R2972 AVDD.n1173 AVDD.t1244 1.4705
R2973 AVDD.n1860 AVDD.n1859 1.46537
R2974 AVDD.n1864 AVDD.n1863 1.46537
R2975 AVDD.n1833 AVDD.n1832 1.46537
R2976 AVDD.n1918 AVDD.n1917 1.46537
R2977 AVDD.n1916 AVDD.n1915 1.46537
R2978 AVDD.n1911 AVDD.n1910 1.46537
R2979 AVDD.n1542 AVDD.n1541 1.46537
R2980 AVDD.n1540 AVDD.n1539 1.46537
R2981 AVDD.n1491 AVDD.n1490 1.46537
R2982 AVDD.n1582 AVDD.n1581 1.46537
R2983 AVDD.n1586 AVDD.n1585 1.46537
R2984 AVDD.n1580 AVDD.n1579 1.46537
R2985 AVDD.n1721 AVDD.n1720 1.46537
R2986 AVDD.n1725 AVDD.n1724 1.46537
R2987 AVDD.n1729 AVDD.n1728 1.46537
R2988 AVDD.n1734 AVDD.n1733 1.46537
R2989 AVDD.n1738 AVDD.n1737 1.46537
R2990 AVDD.n1742 AVDD.n1741 1.46537
R2991 AVDD.n1746 AVDD.n1745 1.46537
R2992 AVDD.n1688 AVDD.n1687 1.46537
R2993 AVDD.n1692 AVDD.n1691 1.46537
R2994 AVDD.n1696 AVDD.n1695 1.46537
R2995 AVDD.n1681 AVDD.n1680 1.46537
R2996 AVDD.n1677 AVDD.n1676 1.46537
R2997 AVDD.n1673 AVDD.n1672 1.46537
R2998 AVDD.n1669 AVDD.n1668 1.46537
R2999 AVDD.n278 AVDD.n277 1.46537
R3000 AVDD.n282 AVDD.n281 1.46537
R3001 AVDD.n286 AVDD.n285 1.46537
R3002 AVDD.n271 AVDD.n270 1.46537
R3003 AVDD.n267 AVDD.n266 1.46537
R3004 AVDD.n263 AVDD.n262 1.46537
R3005 AVDD.n259 AVDD.n258 1.46537
R3006 AVDD.n186 AVDD.n185 1.46537
R3007 AVDD.n190 AVDD.n189 1.46537
R3008 AVDD.n194 AVDD.n193 1.46537
R3009 AVDD.n217 AVDD.n216 1.46537
R3010 AVDD.n221 AVDD.n220 1.46537
R3011 AVDD.n225 AVDD.n224 1.46537
R3012 AVDD.n229 AVDD.n228 1.46537
R3013 AVDD.n1106 AVDD.n1105 1.30325
R3014 AVDD.n1084 AVDD.n1083 1.30325
R3015 AVDD.n1035 AVDD.n1034 1.30325
R3016 AVDD.n1134 AVDD.n1132 1.27338
R3017 AVDD.n1127 AVDD.n1125 1.27338
R3018 AVDD.n1130 AVDD.n1129 1.27228
R3019 AVDD.n957 AVDD.n955 1.27228
R3020 AVDD.n953 AVDD.n951 1.27228
R3021 AVDD.n950 AVDD.n948 1.27228
R3022 AVDD.n53 AVDD.n51 1.27228
R3023 AVDD.n1928 AVDD.n1926 1.27228
R3024 AVDD.n1924 AVDD.n1922 1.27228
R3025 AVDD.n1873 AVDD.n1871 1.27228
R3026 AVDD.n1881 AVDD.n1879 1.27228
R3027 AVDD.n1877 AVDD.n1875 1.27228
R3028 AVDD.n1918 AVDD.n1916 1.27228
R3029 AVDD.n1864 AVDD.n1860 1.27228
R3030 AVDD.n1746 AVDD.n1742 1.27228
R3031 AVDD.n1738 AVDD.n1734 1.27228
R3032 AVDD.n1729 AVDD.n1725 1.27228
R3033 AVDD.n1673 AVDD.n1669 1.27228
R3034 AVDD.n1681 AVDD.n1677 1.27228
R3035 AVDD.n1696 AVDD.n1692 1.27228
R3036 AVDD.n1751 AVDD.n1750 1.27228
R3037 AVDD.n1701 AVDD.n1700 1.27228
R3038 AVDD.n76 AVDD.n74 1.27228
R3039 AVDD.n1594 AVDD.n1592 1.27228
R3040 AVDD.n1598 AVDD.n1596 1.27228
R3041 AVDD.n1550 AVDD.n1548 1.27228
R3042 AVDD.n1555 AVDD.n1553 1.27228
R3043 AVDD.n1559 AVDD.n1557 1.27228
R3044 AVDD.n1586 AVDD.n1582 1.27228
R3045 AVDD.n1542 AVDD.n1540 1.27228
R3046 AVDD.n263 AVDD.n259 1.27228
R3047 AVDD.n271 AVDD.n267 1.27228
R3048 AVDD.n286 AVDD.n282 1.27228
R3049 AVDD.n229 AVDD.n225 1.27228
R3050 AVDD.n221 AVDD.n217 1.27228
R3051 AVDD.n194 AVDD.n190 1.27228
R3052 AVDD.n293 AVDD.n291 1.27228
R3053 AVDD.n236 AVDD.n234 1.27228
R3054 AVDD.n1435 AVDD.t88 1.1382
R3055 AVDD.n1394 AVDD.t175 1.1382
R3056 AVDD.n1977 AVDD.t98 1.1382
R3057 AVDD.n1056 AVDD.t186 1.1382
R3058 AVDD.n1932 AVDD.n1931 1.13692
R3059 AVDD.n1784 AVDD.n54 1.13692
R3060 AVDD.n1601 AVDD.n1600 1.13692
R3061 AVDD.n1453 AVDD.n77 1.13692
R3062 AVDD.n1804 AVDD.n1803 0.9995
R3063 AVDD.n1891 AVDD.n1890 0.9995
R3064 AVDD.n1901 AVDD.n1900 0.9995
R3065 AVDD.n1823 AVDD.n1822 0.9995
R3066 AVDD.n1843 AVDD.n1842 0.9995
R3067 AVDD.n1853 AVDD.n1852 0.9995
R3068 AVDD.n1469 AVDD.n1468 0.9995
R3069 AVDD.n1571 AVDD.n1570 0.9995
R3070 AVDD.n1565 AVDD.n1564 0.9995
R3071 AVDD.n1506 AVDD.n1505 0.9995
R3072 AVDD.n1531 AVDD.n1530 0.9995
R3073 AVDD.n1525 AVDD.n1524 0.9995
R3074 AVDD.n1115 AVDD.n1114 0.9995
R3075 AVDD.n1109 AVDD.n1108 0.9995
R3076 AVDD.n1103 AVDD.n1102 0.9995
R3077 AVDD.n1068 AVDD.n1067 0.9995
R3078 AVDD.n1078 AVDD.n1077 0.9995
R3079 AVDD.n1090 AVDD.n1089 0.9995
R3080 AVDD.n1044 AVDD.n1043 0.9995
R3081 AVDD.n1038 AVDD.n1037 0.9995
R3082 AVDD.n1032 AVDD.n1031 0.9995
R3083 AVDD.n1711 AVDD.n1710 0.991625
R3084 AVDD.n1662 AVDD.n1661 0.991625
R3085 AVDD.n243 AVDD.n242 0.991625
R3086 AVDD.n200 AVDD.n199 0.991625
R3087 AVDD.n1931 AVDD.n1930 0.983405
R3088 AVDD.n1920 AVDD.n1784 0.983405
R3089 AVDD.n1600 AVDD.n1599 0.983405
R3090 AVDD.n1589 AVDD.n1453 0.983405
R3091 AVDD.n1132 AVDD.n1130 0.937025
R3092 AVDD.n951 AVDD.n950 0.937025
R3093 AVDD.n1884 AVDD.n1883 0.822966
R3094 AVDD.n1906 AVDD.n1785 0.822966
R3095 AVDD.n1561 AVDD.n1560 0.822966
R3096 AVDD.n1575 AVDD.n1454 0.822966
R3097 AVDD.n1748 AVDD.n1747 0.737223
R3098 AVDD.n1665 AVDD.n1635 0.737223
R3099 AVDD.n1755 AVDD.n63 0.737223
R3100 AVDD.n1705 AVDD.n1698 0.737223
R3101 AVDD.n289 AVDD.n288 0.737223
R3102 AVDD.n212 AVDD.n176 0.737223
R3103 AVDD.n294 AVDD.n143 0.737223
R3104 AVDD.n237 AVDD.n230 0.737223
R3105 AVDD.n1714 AVDD.n1635 0.725061
R3106 AVDD.n1706 AVDD.n1705 0.725061
R3107 AVDD.n255 AVDD.n176 0.725061
R3108 AVDD.n238 AVDD.n237 0.725061
R3109 AVDD.n1112 AVDD.n1111 0.66425
R3110 AVDD.n1074 AVDD.n1073 0.66425
R3111 AVDD.n1041 AVDD.n1040 0.66425
R3112 AVDD.n1930 AVDD.n46 0.639318
R3113 AVDD.n1883 AVDD.n1866 0.639318
R3114 AVDD.n1920 AVDD.n1919 0.639318
R3115 AVDD.n1858 AVDD.n1785 0.639318
R3116 AVDD.n1599 AVDD.n69 0.639318
R3117 AVDD.n1560 AVDD.n1543 0.639318
R3118 AVDD.n1589 AVDD.n1588 0.639318
R3119 AVDD.n1535 AVDD.n1454 0.639318
R3120 AVDD.n1884 AVDD.n46 0.585196
R3121 AVDD.n1919 AVDD.n1906 0.585196
R3122 AVDD.n1747 AVDD.n1714 0.585196
R3123 AVDD.n1706 AVDD.n63 0.585196
R3124 AVDD.n1561 AVDD.n69 0.585196
R3125 AVDD.n1588 AVDD.n1575 0.585196
R3126 AVDD.n288 AVDD.n255 0.585196
R3127 AVDD.n238 AVDD.n143 0.585196
R3128 AVDD.n1929 AVDD.n53 0.236091
R3129 AVDD.n1882 AVDD.n1873 0.236091
R3130 AVDD.n1590 AVDD.n76 0.236091
R3131 AVDD.n1551 AVDD.n1550 0.236091
R3132 AVDD.n980 AVDD.n979 0.166289
R3133 AVDD.n1052 AVDD.n1051 0.166289
R3134 AVDD.n1053 AVDD.n1052 0.166289
R3135 AVDD.n1730 AVDD.n1729 0.150184
R3136 AVDD.n1697 AVDD.n1696 0.150184
R3137 AVDD.n287 AVDD.n286 0.150184
R3138 AVDD.n213 AVDD.n194 0.150184
R3139 AVDD.n1794 AVDD.n1792 0.14
R3140 AVDD.n1798 AVDD.n1792 0.14
R3141 AVDD.n1799 AVDD.n1791 0.14
R3142 AVDD.n1803 AVDD.n1791 0.14
R3143 AVDD.n1804 AVDD.n1790 0.14
R3144 AVDD.n1808 AVDD.n1790 0.14
R3145 AVDD.n1886 AVDD.n1789 0.14
R3146 AVDD.n1890 AVDD.n1789 0.14
R3147 AVDD.n1891 AVDD.n1788 0.14
R3148 AVDD.n1895 AVDD.n1788 0.14
R3149 AVDD.n1896 AVDD.n1787 0.14
R3150 AVDD.n1900 AVDD.n1787 0.14
R3151 AVDD.n1901 AVDD.n1786 0.14
R3152 AVDD.n1905 AVDD.n1786 0.14
R3153 AVDD.n1813 AVDD.n1811 0.14
R3154 AVDD.n1817 AVDD.n1811 0.14
R3155 AVDD.n1818 AVDD.n1810 0.14
R3156 AVDD.n1822 AVDD.n1810 0.14
R3157 AVDD.n1823 AVDD.n1809 0.14
R3158 AVDD.n1827 AVDD.n1809 0.14
R3159 AVDD.n1838 AVDD.n1837 0.14
R3160 AVDD.n1842 AVDD.n1837 0.14
R3161 AVDD.n1843 AVDD.n1836 0.14
R3162 AVDD.n1847 AVDD.n1836 0.14
R3163 AVDD.n1848 AVDD.n1835 0.14
R3164 AVDD.n1852 AVDD.n1835 0.14
R3165 AVDD.n1853 AVDD.n1834 0.14
R3166 AVDD.n1857 AVDD.n1834 0.14
R3167 AVDD.n1713 AVDD.n1636 0.14
R3168 AVDD.n1711 AVDD.n1636 0.14
R3169 AVDD.n1710 AVDD.n1638 0.14
R3170 AVDD.n1708 AVDD.n1638 0.14
R3171 AVDD.n1646 AVDD.n1641 0.14
R3172 AVDD.n1644 AVDD.n1641 0.14
R3173 AVDD.n1664 AVDD.n1654 0.14
R3174 AVDD.n1662 AVDD.n1654 0.14
R3175 AVDD.n1661 AVDD.n1656 0.14
R3176 AVDD.n1659 AVDD.n1656 0.14
R3177 AVDD.n1652 AVDD.n1647 0.14
R3178 AVDD.n1650 AVDD.n1647 0.14
R3179 AVDD.n1459 AVDD.n1457 0.14
R3180 AVDD.n1463 AVDD.n1457 0.14
R3181 AVDD.n1464 AVDD.n1456 0.14
R3182 AVDD.n1468 AVDD.n1456 0.14
R3183 AVDD.n1469 AVDD.n1455 0.14
R3184 AVDD.n1473 AVDD.n1455 0.14
R3185 AVDD.n1573 AVDD.n1474 0.14
R3186 AVDD.n1571 AVDD.n1474 0.14
R3187 AVDD.n1570 AVDD.n1477 0.14
R3188 AVDD.n1568 AVDD.n1477 0.14
R3189 AVDD.n1567 AVDD.n1480 0.14
R3190 AVDD.n1565 AVDD.n1480 0.14
R3191 AVDD.n1564 AVDD.n1483 0.14
R3192 AVDD.n1562 AVDD.n1483 0.14
R3193 AVDD.n1496 AVDD.n1494 0.14
R3194 AVDD.n1500 AVDD.n1494 0.14
R3195 AVDD.n1501 AVDD.n1493 0.14
R3196 AVDD.n1505 AVDD.n1493 0.14
R3197 AVDD.n1506 AVDD.n1492 0.14
R3198 AVDD.n1510 AVDD.n1492 0.14
R3199 AVDD.n1533 AVDD.n1511 0.14
R3200 AVDD.n1531 AVDD.n1511 0.14
R3201 AVDD.n1530 AVDD.n1514 0.14
R3202 AVDD.n1528 AVDD.n1514 0.14
R3203 AVDD.n1527 AVDD.n1517 0.14
R3204 AVDD.n1525 AVDD.n1517 0.14
R3205 AVDD.n1524 AVDD.n1520 0.14
R3206 AVDD.n1520 AVDD.n1486 0.14
R3207 AVDD.n239 AVDD.n178 0.14
R3208 AVDD.n242 AVDD.n178 0.14
R3209 AVDD.n243 AVDD.n177 0.14
R3210 AVDD.n247 AVDD.n177 0.14
R3211 AVDD.n253 AVDD.n248 0.14
R3212 AVDD.n251 AVDD.n248 0.14
R3213 AVDD.n196 AVDD.n179 0.14
R3214 AVDD.n199 AVDD.n196 0.14
R3215 AVDD.n200 AVDD.n195 0.14
R3216 AVDD.n204 AVDD.n195 0.14
R3217 AVDD.n210 AVDD.n205 0.14
R3218 AVDD.n208 AVDD.n205 0.14
R3219 AVDD.n1117 AVDD.n666 0.14
R3220 AVDD.n1115 AVDD.n666 0.14
R3221 AVDD.n1114 AVDD.n669 0.14
R3222 AVDD.n1112 AVDD.n669 0.14
R3223 AVDD.n1111 AVDD.n672 0.14
R3224 AVDD.n1109 AVDD.n672 0.14
R3225 AVDD.n1108 AVDD.n674 0.14
R3226 AVDD.n1106 AVDD.n674 0.14
R3227 AVDD.n1105 AVDD.n677 0.14
R3228 AVDD.n1103 AVDD.n677 0.14
R3229 AVDD.n1102 AVDD.n680 0.14
R3230 AVDD.n1100 AVDD.n680 0.14
R3231 AVDD.n1062 AVDD.n692 0.14
R3232 AVDD.n1067 AVDD.n692 0.14
R3233 AVDD.n1068 AVDD.n691 0.14
R3234 AVDD.n1073 AVDD.n691 0.14
R3235 AVDD.n1074 AVDD.n690 0.14
R3236 AVDD.n1077 AVDD.n690 0.14
R3237 AVDD.n1078 AVDD.n689 0.14
R3238 AVDD.n1083 AVDD.n689 0.14
R3239 AVDD.n1084 AVDD.n688 0.14
R3240 AVDD.n1089 AVDD.n688 0.14
R3241 AVDD.n1090 AVDD.n687 0.14
R3242 AVDD.n1095 AVDD.n687 0.14
R3243 AVDD.n1046 AVDD.n901 0.14
R3244 AVDD.n1044 AVDD.n901 0.14
R3245 AVDD.n1043 AVDD.n904 0.14
R3246 AVDD.n1041 AVDD.n904 0.14
R3247 AVDD.n1040 AVDD.n907 0.14
R3248 AVDD.n1038 AVDD.n907 0.14
R3249 AVDD.n1037 AVDD.n909 0.14
R3250 AVDD.n1035 AVDD.n909 0.14
R3251 AVDD.n1034 AVDD.n912 0.14
R3252 AVDD.n1032 AVDD.n912 0.14
R3253 AVDD.n1031 AVDD.n915 0.14
R3254 AVDD.n1029 AVDD.n915 0.14
R3255 AVDD.n933 AVDD.n897 0.13175
R3256 AVDD.n978 AVDD.n897 0.13175
R3257 AVDD.n930 AVDD.n898 0.13175
R3258 AVDD.n978 AVDD.n898 0.13175
R3259 AVDD.n1156 AVDD.n1155 0.105779
R3260 AVDD.n1149 AVDD.n1148 0.105779
R3261 AVDD.n312 AVDD.n311 0.103153
R3262 AVDD.n548 AVDD.n547 0.103153
R3263 AVDD.n1213 AVDD.n1212 0.101802
R3264 AVDD.n750 AVDD.n746 0.101802
R3265 AVDD.n1212 AVDD.n1211 0.101802
R3266 AVDD.n1226 AVDD.n653 0.101802
R3267 AVDD.n1226 AVDD.n1225 0.101802
R3268 AVDD.n750 AVDD.n749 0.101802
R3269 AVDD.n1885 AVDD.n1808 0.10175
R3270 AVDD.n1828 AVDD.n1827 0.10175
R3271 AVDD.n1574 AVDD.n1473 0.10175
R3272 AVDD.n1534 AVDD.n1510 0.10175
R3273 AVDD.n344 AVDD.n321 0.0992755
R3274 AVDD.n345 AVDD.n344 0.0992755
R3275 AVDD.n562 AVDD.n354 0.0992755
R3276 AVDD.n562 AVDD.n561 0.0992755
R3277 AVDD.n469 AVDD.n465 0.0992755
R3278 AVDD.n469 AVDD.n468 0.0992755
R3279 AVDD.n554 AVDD.n553 0.0931471
R3280 AVDD.n555 AVDD.n554 0.0931471
R3281 AVDD.n510 AVDD.n509 0.0931471
R3282 AVDD.n509 AVDD.n106 0.0931471
R3283 AVDD.n510 AVDD.n107 0.0931471
R3284 AVDD.n1409 AVDD.n107 0.0931471
R3285 AVDD.n840 AVDD.n20 0.0931471
R3286 AVDD.n37 AVDD.n20 0.0931471
R3287 AVDD.n840 AVDD.n38 0.0931471
R3288 AVDD.n1951 AVDD.n38 0.0931471
R3289 AVDD.n1154 AVDD.n1153 0.0931471
R3290 AVDD.n1219 AVDD.n1154 0.0931471
R3291 AVDD.n557 AVDD.n556 0.0931471
R3292 AVDD.n556 AVDD.n555 0.0931471
R3293 AVDD.n442 AVDD.n441 0.0931471
R3294 AVDD.n441 AVDD.n106 0.0931471
R3295 AVDD.n442 AVDD.n108 0.0931471
R3296 AVDD.n1409 AVDD.n108 0.0931471
R3297 AVDD.n826 AVDD.n825 0.0931471
R3298 AVDD.n825 AVDD.n37 0.0931471
R3299 AVDD.n826 AVDD.n39 0.0931471
R3300 AVDD.n1951 AVDD.n39 0.0931471
R3301 AVDD.n349 AVDD.n91 0.0931471
R3302 AVDD.n555 AVDD.n91 0.0931471
R3303 AVDD.n1411 AVDD.n92 0.0931471
R3304 AVDD.n106 AVDD.n92 0.0931471
R3305 AVDD.n1411 AVDD.n1410 0.0931471
R3306 AVDD.n1410 AVDD.n1409 0.0931471
R3307 AVDD.n317 AVDD.n83 0.0931471
R3308 AVDD.n555 AVDD.n83 0.0931471
R3309 AVDD.n1407 AVDD.n84 0.0931471
R3310 AVDD.n106 AVDD.n84 0.0931471
R3311 AVDD.n1408 AVDD.n1407 0.0931471
R3312 AVDD.n1409 AVDD.n1408 0.0931471
R3313 AVDD.n1218 AVDD.n1217 0.0931471
R3314 AVDD.n1219 AVDD.n1218 0.0931471
R3315 AVDD.n1207 AVDD.n656 0.0931471
R3316 AVDD.n1219 AVDD.n656 0.0931471
R3317 AVDD.n1221 AVDD.n1220 0.0931471
R3318 AVDD.n1220 AVDD.n1219 0.0931471
R3319 AVDD.n1953 AVDD.n23 0.0931471
R3320 AVDD.n37 AVDD.n23 0.0931471
R3321 AVDD.n1953 AVDD.n1952 0.0931471
R3322 AVDD.n1952 AVDD.n1951 0.0931471
R3323 AVDD.n1949 AVDD.n1943 0.0931471
R3324 AVDD.n1943 AVDD.n37 0.0931471
R3325 AVDD.n1950 AVDD.n1949 0.0931471
R3326 AVDD.n1951 AVDD.n1950 0.0931471
R3327 AVDD.n2000 AVDD.n14 0.0931471
R3328 AVDD.n14 AVDD.n5 0.0931471
R3329 AVDD.n2000 AVDD.n7 0.0931471
R3330 AVDD.n2016 AVDD.n7 0.0931471
R3331 AVDD.n2014 AVDD.n11 0.0931471
R3332 AVDD.n11 AVDD.n5 0.0931471
R3333 AVDD.n2015 AVDD.n2014 0.0931471
R3334 AVDD.n2016 AVDD.n2015 0.0931471
R3335 AVDD.n1365 AVDD.n1364 0.0931471
R3336 AVDD.n1364 AVDD.n5 0.0931471
R3337 AVDD.n1365 AVDD.n6 0.0931471
R3338 AVDD.n2016 AVDD.n6 0.0931471
R3339 AVDD.n2018 AVDD.n1 0.0931471
R3340 AVDD.n5 AVDD.n1 0.0931471
R3341 AVDD.n2018 AVDD.n2017 0.0931471
R3342 AVDD.n2017 AVDD.n2016 0.0931471
R3343 AVDD.n1060 AVDD.n1059 0.0737558
R3344 AVDD.n1059 AVDD.n1058 0.0737558
R3345 AVDD.n1054 AVDD.n686 0.0737558
R3346 AVDD.n1217 AVDD.n1216 0.0723953
R3347 AVDD.n1153 AVDD.n1152 0.0723953
R3348 AVDD.n1207 AVDD.n1206 0.0723953
R3349 AVDD.n1221 AVDD.n654 0.0723953
R3350 AVDD.n989 AVDD.n987 0.0720299
R3351 AVDD.n318 AVDD.n317 0.070602
R3352 AVDD.n1028 AVDD.n1027 0.0692176
R3353 AVDD.n895 AVDD.n894 0.0682419
R3354 AVDD.n1055 AVDD.n895 0.0682419
R3355 AVDD.n1011 AVDD.n896 0.0682419
R3356 AVDD.n1055 AVDD.n896 0.0682419
R3357 AVDD.n456 AVDD.n89 0.0682419
R3358 AVDD.n1435 AVDD.n89 0.0682419
R3359 AVDD.n424 AVDD.n113 0.0682419
R3360 AVDD.n1394 AVDD.n113 0.0682419
R3361 AVDD.n788 AVDD.n22 0.0682419
R3362 AVDD.n1977 AVDD.n22 0.0682419
R3363 AVDD.n767 AVDD.n657 0.0682419
R3364 AVDD.n1056 AVDD.n657 0.0682419
R3365 AVDD.n134 AVDD.n90 0.0682419
R3366 AVDD.n1435 AVDD.n90 0.0682419
R3367 AVDD.n1393 AVDD.n1392 0.0682419
R3368 AVDD.n1394 AVDD.n1393 0.0682419
R3369 AVDD.n1434 AVDD.n1433 0.0682419
R3370 AVDD.n1435 AVDD.n1434 0.0682419
R3371 AVDD.n110 AVDD.n104 0.0682419
R3372 AVDD.n1394 AVDD.n104 0.0682419
R3373 AVDD.n1976 AVDD.n1975 0.0682419
R3374 AVDD.n1977 AVDD.n1976 0.0682419
R3375 AVDD.n1437 AVDD.n1436 0.0682419
R3376 AVDD.n1436 AVDD.n1435 0.0682419
R3377 AVDD.n1768 AVDD.n40 0.0682419
R3378 AVDD.n1056 AVDD.n40 0.0682419
R3379 AVDD.n1168 AVDD.n35 0.0682419
R3380 AVDD.n1056 AVDD.n35 0.0682419
R3381 AVDD.n1279 AVDD.n8 0.0682419
R3382 AVDD.n1977 AVDD.n8 0.0682419
R3383 AVDD.n1243 AVDD.n644 0.0682419
R3384 AVDD.n1056 AVDD.n644 0.0682419
R3385 AVDD.n1622 AVDD.n3 0.0682419
R3386 AVDD.n1977 AVDD.n3 0.0682419
R3387 AVDD.n163 AVDD.n109 0.0682419
R3388 AVDD.n1394 AVDD.n109 0.0682419
R3389 AVDD.n532 AVDD.n88 0.0668158
R3390 AVDD.n1435 AVDD.n88 0.0668158
R3391 AVDD.n383 AVDD.n112 0.0668158
R3392 AVDD.n1394 AVDD.n112 0.0668158
R3393 AVDD.n1979 AVDD.n1978 0.0668158
R3394 AVDD.n1978 AVDD.n1977 0.0668158
R3395 AVDD.n704 AVDD.n658 0.0668158
R3396 AVDD.n1056 AVDD.n658 0.0668158
R3397 AVDD.n456 AVDD.n87 0.0668158
R3398 AVDD.n1435 AVDD.n87 0.0668158
R3399 AVDD.n424 AVDD.n111 0.0668158
R3400 AVDD.n1394 AVDD.n111 0.0668158
R3401 AVDD.n788 AVDD.n9 0.0668158
R3402 AVDD.n1977 AVDD.n9 0.0668158
R3403 AVDD.n767 AVDD.n655 0.0668158
R3404 AVDD.n1056 AVDD.n655 0.0668158
R3405 AVDD.n134 AVDD.n86 0.0668158
R3406 AVDD.n1435 AVDD.n86 0.0668158
R3407 AVDD.n1392 AVDD.n105 0.0668158
R3408 AVDD.n1394 AVDD.n105 0.0668158
R3409 AVDD.n1433 AVDD.n85 0.0668158
R3410 AVDD.n1435 AVDD.n85 0.0668158
R3411 AVDD.n1395 AVDD.n110 0.0668158
R3412 AVDD.n1395 AVDD.n1394 0.0668158
R3413 AVDD.n1975 AVDD.n4 0.0668158
R3414 AVDD.n1977 AVDD.n4 0.0668158
R3415 AVDD.n1168 AVDD.n41 0.0668158
R3416 AVDD.n1056 AVDD.n41 0.0668158
R3417 AVDD.n1279 AVDD.n21 0.0668158
R3418 AVDD.n1977 AVDD.n21 0.0668158
R3419 AVDD.n1243 AVDD.n36 0.0668158
R3420 AVDD.n1056 AVDD.n36 0.0668158
R3421 AVDD.n351 AVDD.n350 0.0660102
R3422 AVDD.n462 AVDD.n355 0.0660102
R3423 AVDD.n1217 AVDD.n1159 0.0629767
R3424 AVDD.n1153 AVDD.n659 0.0629767
R3425 AVDD.n1208 AVDD.n1207 0.0629767
R3426 AVDD.n1222 AVDD.n1221 0.0629767
R3427 AVDD.n1137 AVDD.n1135 0.0619118
R3428 AVDD.n1123 AVDD.n664 0.0616241
R3429 AVDD.n349 AVDD.n348 0.0614184
R3430 AVDD.n558 AVDD.n557 0.0614184
R3431 AVDD.n553 AVDD.n356 0.0614184
R3432 AVDD.n1398 AVDD.n1397 0.0525345
R3433 AVDD.n1403 AVDD.n1402 0.0525345
R3434 AVDD.n1416 AVDD.n1415 0.0525345
R3435 AVDD.n447 AVDD.n446 0.0525345
R3436 AVDD.n505 AVDD.n504 0.0525345
R3437 AVDD.n515 AVDD.n514 0.0525345
R3438 AVDD.n831 AVDD.n830 0.0525345
R3439 AVDD.n836 AVDD.n835 0.0525345
R3440 AVDD.n1939 AVDD.n1938 0.0525345
R3441 AVDD.n1945 AVDD.n1944 0.0525345
R3442 AVDD.n1958 AVDD.n1957 0.0525345
R3443 AVDD.n989 AVDD.n988 0.0513315
R3444 AVDD.n941 AVDD.n686 0.0507941
R3445 AVDD.n597 AVDD.n124 0.050569
R3446 AVDD.n597 AVDD.n125 0.050569
R3447 AVDD.n1262 AVDD.n635 0.050569
R3448 AVDD.n845 AVDD.n844 0.050569
R3449 AVDD.n1262 AVDD.n1261 0.050569
R3450 AVDD.n996 AVDD.n995 0.0465048
R3451 AVDD.n974 AVDD.n973 0.0445515
R3452 AVDD.n963 AVDD.n962 0.0440678
R3453 AVDD.n992 AVDD.n991 0.0436757
R3454 AVDD.n993 AVDD.n992 0.0436757
R3455 AVDD.n993 AVDD.n929 0.0436757
R3456 AVDD.n995 AVDD.n929 0.0436757
R3457 AVDD.n971 AVDD.n931 0.0433141
R3458 AVDD.n970 AVDD.n931 0.0433141
R3459 AVDD.n969 AVDD.n932 0.0433141
R3460 AVDD.n967 AVDD.n966 0.0433141
R3461 AVDD.n966 AVDD.n965 0.0433141
R3462 AVDD.n965 AVDD.n934 0.0433141
R3463 AVDD.n963 AVDD.n934 0.0433141
R3464 AVDD.n972 AVDD.n971 0.0430669
R3465 AVDD.n1097 AVDD.n1096 0.0430647
R3466 AVDD.n1061 AVDD.n693 0.0428653
R3467 AVDD.n684 AVDD.n683 0.0417941
R3468 AVDD.n944 AVDD.n943 0.0417941
R3469 AVDD.n552 AVDD.n551 0.0417245
R3470 AVDD.n1121 AVDD.n1120 0.0416007
R3471 AVDD.n1135 AVDD.n663 0.0415824
R3472 AVDD.n1123 AVDD.n1122 0.0413899
R3473 AVDD.n1158 AVDD.n1157 0.041314
R3474 AVDD.n1215 AVDD.n1214 0.041314
R3475 AVDD.n745 AVDD.n744 0.041314
R3476 AVDD.n1151 AVDD.n1150 0.041314
R3477 AVDD.n1210 AVDD.n1209 0.041314
R3478 AVDD.n1205 AVDD.n1204 0.041314
R3479 AVDD.n1224 AVDD.n1223 0.041314
R3480 AVDD.n748 AVDD.n747 0.041314
R3481 AVDD.n970 AVDD.n969 0.040902
R3482 AVDD.n314 AVDD.n313 0.0402959
R3483 AVDD.n320 AVDD.n319 0.0402959
R3484 AVDD.n347 AVDD.n346 0.0402959
R3485 AVDD.n353 AVDD.n352 0.0402959
R3486 AVDD.n560 AVDD.n559 0.0402959
R3487 AVDD.n464 AVDD.n463 0.0402959
R3488 AVDD.n467 AVDD.n466 0.0402959
R3489 AVDD.n550 AVDD.n549 0.0402959
R3490 AVDD.n1147 AVDD.n1146 0.0395167
R3491 AVDD.n1026 AVDD.n1025 0.0394276
R3492 AVDD.n546 AVDD.n545 0.0393731
R3493 AVDD.n1782 AVDD.n56 0.0392688
R3494 AVDD.n310 AVDD.n309 0.0391565
R3495 AVDD.n946 AVDD.n945 0.0387235
R3496 AVDD.n1028 AVDD.n918 0.0383
R3497 AVDD.n946 AVDD.n942 0.0373471
R3498 AVDD.n1099 AVDD.n1098 0.0371353
R3499 AVDD.n1118 AVDD.n665 0.0369637
R3500 AVDD.n1099 AVDD.n685 0.0369235
R3501 AVDD.n1119 AVDD.n1118 0.0367529
R3502 AVDD.n1407 AVDD.n1406 0.0360345
R3503 AVDD.n1411 AVDD.n103 0.0360345
R3504 AVDD.n443 AVDD.n442 0.0360345
R3505 AVDD.n511 AVDD.n510 0.0360345
R3506 AVDD.n827 AVDD.n826 0.0360345
R3507 AVDD.n841 AVDD.n840 0.0360345
R3508 AVDD.n1949 AVDD.n1948 0.0360345
R3509 AVDD.n1953 AVDD.n34 0.0360345
R3510 AVDD.n1060 AVDD.n694 0.0359624
R3511 AVDD.n1936 AVDD.n42 0.0347688
R3512 AVDD.n1451 AVDD.n79 0.0347688
R3513 AVDD.n998 AVDD.n997 0.0347688
R3514 AVDD.n1607 AVDD.n1606 0.0347688
R3515 AVDD.n1936 AVDD.n1935 0.0347688
R3516 AVDD.n148 AVDD.n79 0.0347688
R3517 AVDD.n1606 AVDD.n1604 0.0347688
R3518 AVDD.n317 AVDD.n316 0.0345816
R3519 AVDD.n62 AVDD.n42 0.0341759
R3520 AVDD.n1757 AVDD.n61 0.0341759
R3521 AVDD.n1760 AVDD.n61 0.0341759
R3522 AVDD.n1761 AVDD.n1760 0.0341759
R3523 AVDD.n1762 AVDD.n1761 0.0341759
R3524 AVDD.n1762 AVDD.n60 0.0341759
R3525 AVDD.n1764 AVDD.n60 0.0341759
R3526 AVDD.n1765 AVDD.n59 0.0341759
R3527 AVDD.n1767 AVDD.n59 0.0341759
R3528 AVDD.n1770 AVDD.n1769 0.0341759
R3529 AVDD.n1770 AVDD.n58 0.0341759
R3530 AVDD.n1772 AVDD.n58 0.0341759
R3531 AVDD.n1774 AVDD.n1773 0.0341759
R3532 AVDD.n1775 AVDD.n1774 0.0341759
R3533 AVDD.n1775 AVDD.n57 0.0341759
R3534 AVDD.n1778 AVDD.n57 0.0341759
R3535 AVDD.n1779 AVDD.n1778 0.0341759
R3536 AVDD.n1780 AVDD.n1779 0.0341759
R3537 AVDD.n309 AVDD.n142 0.0341759
R3538 AVDD.n307 AVDD.n306 0.0341759
R3539 AVDD.n306 AVDD.n305 0.0341759
R3540 AVDD.n305 AVDD.n296 0.0341759
R3541 AVDD.n302 AVDD.n296 0.0341759
R3542 AVDD.n302 AVDD.n301 0.0341759
R3543 AVDD.n301 AVDD.n300 0.0341759
R3544 AVDD.n299 AVDD.n297 0.0341759
R3545 AVDD.n297 AVDD.n82 0.0341759
R3546 AVDD.n1439 AVDD.n1438 0.0341759
R3547 AVDD.n1439 AVDD.n81 0.0341759
R3548 AVDD.n1441 AVDD.n81 0.0341759
R3549 AVDD.n1443 AVDD.n1442 0.0341759
R3550 AVDD.n1444 AVDD.n1443 0.0341759
R3551 AVDD.n1444 AVDD.n80 0.0341759
R3552 AVDD.n1447 AVDD.n80 0.0341759
R3553 AVDD.n1448 AVDD.n1447 0.0341759
R3554 AVDD.n1449 AVDD.n1448 0.0341759
R3555 AVDD.n999 AVDD.n998 0.0341759
R3556 AVDD.n1000 AVDD.n999 0.0341759
R3557 AVDD.n1000 AVDD.n924 0.0341759
R3558 AVDD.n1003 AVDD.n924 0.0341759
R3559 AVDD.n1004 AVDD.n1003 0.0341759
R3560 AVDD.n1005 AVDD.n1004 0.0341759
R3561 AVDD.n1005 AVDD.n923 0.0341759
R3562 AVDD.n1007 AVDD.n923 0.0341759
R3563 AVDD.n1008 AVDD.n922 0.0341759
R3564 AVDD.n1010 AVDD.n922 0.0341759
R3565 AVDD.n1013 AVDD.n1012 0.0341759
R3566 AVDD.n1013 AVDD.n921 0.0341759
R3567 AVDD.n1015 AVDD.n921 0.0341759
R3568 AVDD.n1017 AVDD.n1016 0.0341759
R3569 AVDD.n1018 AVDD.n1017 0.0341759
R3570 AVDD.n1018 AVDD.n920 0.0341759
R3571 AVDD.n1021 AVDD.n920 0.0341759
R3572 AVDD.n1022 AVDD.n1021 0.0341759
R3573 AVDD.n1023 AVDD.n1022 0.0341759
R3574 AVDD.n1023 AVDD.n919 0.0341759
R3575 AVDD.n1025 AVDD.n919 0.0341759
R3576 AVDD.n1607 AVDD.n64 0.0341759
R3577 AVDD.n1633 AVDD.n65 0.0341759
R3578 AVDD.n1630 AVDD.n65 0.0341759
R3579 AVDD.n1630 AVDD.n1629 0.0341759
R3580 AVDD.n1629 AVDD.n1628 0.0341759
R3581 AVDD.n1628 AVDD.n1608 0.0341759
R3582 AVDD.n1626 AVDD.n1608 0.0341759
R3583 AVDD.n1625 AVDD.n1609 0.0341759
R3584 AVDD.n1623 AVDD.n1609 0.0341759
R3585 AVDD.n1621 AVDD.n1620 0.0341759
R3586 AVDD.n1620 AVDD.n1610 0.0341759
R3587 AVDD.n1618 AVDD.n1610 0.0341759
R3588 AVDD.n1617 AVDD.n1611 0.0341759
R3589 AVDD.n1615 AVDD.n1611 0.0341759
R3590 AVDD.n1615 AVDD.n1614 0.0341759
R3591 AVDD.n1614 AVDD.n1613 0.0341759
R3592 AVDD.n1613 AVDD.n44 0.0341759
R3593 AVDD.n1933 AVDD.n44 0.0341759
R3594 AVDD.n148 AVDD.n146 0.0341759
R3595 AVDD.n174 AVDD.n147 0.0341759
R3596 AVDD.n171 AVDD.n147 0.0341759
R3597 AVDD.n171 AVDD.n170 0.0341759
R3598 AVDD.n170 AVDD.n169 0.0341759
R3599 AVDD.n169 AVDD.n149 0.0341759
R3600 AVDD.n167 AVDD.n149 0.0341759
R3601 AVDD.n166 AVDD.n150 0.0341759
R3602 AVDD.n164 AVDD.n150 0.0341759
R3603 AVDD.n162 AVDD.n161 0.0341759
R3604 AVDD.n161 AVDD.n151 0.0341759
R3605 AVDD.n159 AVDD.n151 0.0341759
R3606 AVDD.n158 AVDD.n152 0.0341759
R3607 AVDD.n156 AVDD.n152 0.0341759
R3608 AVDD.n156 AVDD.n155 0.0341759
R3609 AVDD.n155 AVDD.n154 0.0341759
R3610 AVDD.n154 AVDD.n67 0.0341759
R3611 AVDD.n1602 AVDD.n67 0.0341759
R3612 AVDD.n517 AVDD.n396 0.0337609
R3613 AVDD.n1993 AVDD.n15 0.0337609
R3614 AVDD.n518 AVDD.n517 0.0337609
R3615 AVDD.n1993 AVDD.n1992 0.0337609
R3616 AVDD.n396 AVDD.n364 0.0331854
R3617 AVDD.n394 AVDD.n364 0.0331854
R3618 AVDD.n394 AVDD.n393 0.0331854
R3619 AVDD.n393 AVDD.n392 0.0331854
R3620 AVDD.n392 AVDD.n365 0.0331854
R3621 AVDD.n389 AVDD.n365 0.0331854
R3622 AVDD.n389 AVDD.n388 0.0331854
R3623 AVDD.n388 AVDD.n387 0.0331854
R3624 AVDD.n386 AVDD.n366 0.0331854
R3625 AVDD.n384 AVDD.n366 0.0331854
R3626 AVDD.n382 AVDD.n381 0.0331854
R3627 AVDD.n381 AVDD.n367 0.0331854
R3628 AVDD.n379 AVDD.n367 0.0331854
R3629 AVDD.n378 AVDD.n368 0.0331854
R3630 AVDD.n376 AVDD.n368 0.0331854
R3631 AVDD.n376 AVDD.n375 0.0331854
R3632 AVDD.n375 AVDD.n374 0.0331854
R3633 AVDD.n374 AVDD.n369 0.0331854
R3634 AVDD.n371 AVDD.n369 0.0331854
R3635 AVDD.n371 AVDD.n370 0.0331854
R3636 AVDD.n370 AVDD.n15 0.0331854
R3637 AVDD.n545 AVDD.n358 0.0331854
R3638 AVDD.n543 AVDD.n358 0.0331854
R3639 AVDD.n543 AVDD.n542 0.0331854
R3640 AVDD.n542 AVDD.n541 0.0331854
R3641 AVDD.n541 AVDD.n359 0.0331854
R3642 AVDD.n538 AVDD.n359 0.0331854
R3643 AVDD.n538 AVDD.n537 0.0331854
R3644 AVDD.n537 AVDD.n536 0.0331854
R3645 AVDD.n535 AVDD.n360 0.0331854
R3646 AVDD.n533 AVDD.n360 0.0331854
R3647 AVDD.n531 AVDD.n530 0.0331854
R3648 AVDD.n530 AVDD.n361 0.0331854
R3649 AVDD.n528 AVDD.n361 0.0331854
R3650 AVDD.n527 AVDD.n362 0.0331854
R3651 AVDD.n525 AVDD.n362 0.0331854
R3652 AVDD.n525 AVDD.n524 0.0331854
R3653 AVDD.n524 AVDD.n523 0.0331854
R3654 AVDD.n523 AVDD.n363 0.0331854
R3655 AVDD.n520 AVDD.n363 0.0331854
R3656 AVDD.n520 AVDD.n519 0.0331854
R3657 AVDD.n519 AVDD.n518 0.0331854
R3658 AVDD.n1144 AVDD.n1143 0.0331854
R3659 AVDD.n1144 AVDD.n660 0.0331854
R3660 AVDD.n1146 AVDD.n660 0.0331854
R3661 AVDD.n1992 AVDD.n16 0.0331854
R3662 AVDD.n1990 AVDD.n16 0.0331854
R3663 AVDD.n1990 AVDD.n1989 0.0331854
R3664 AVDD.n1989 AVDD.n1988 0.0331854
R3665 AVDD.n1988 AVDD.n17 0.0331854
R3666 AVDD.n1985 AVDD.n17 0.0331854
R3667 AVDD.n1985 AVDD.n1984 0.0331854
R3668 AVDD.n1984 AVDD.n1983 0.0331854
R3669 AVDD.n1982 AVDD.n18 0.0331854
R3670 AVDD.n1980 AVDD.n18 0.0331854
R3671 AVDD.n851 AVDD.n19 0.0331854
R3672 AVDD.n851 AVDD.n850 0.0331854
R3673 AVDD.n853 AVDD.n850 0.0331854
R3674 AVDD.n854 AVDD.n849 0.0331854
R3675 AVDD.n856 AVDD.n849 0.0331854
R3676 AVDD.n857 AVDD.n856 0.0331854
R3677 AVDD.n860 AVDD.n857 0.0331854
R3678 AVDD.n1765 AVDD.n1764 0.0325158
R3679 AVDD.n1773 AVDD.n1772 0.0325158
R3680 AVDD.n300 AVDD.n299 0.0325158
R3681 AVDD.n1442 AVDD.n1441 0.0325158
R3682 AVDD.n1008 AVDD.n1007 0.0325158
R3683 AVDD.n1016 AVDD.n1015 0.0325158
R3684 AVDD.n1626 AVDD.n1625 0.0325158
R3685 AVDD.n1618 AVDD.n1617 0.0325158
R3686 AVDD.n167 AVDD.n166 0.0325158
R3687 AVDD.n159 AVDD.n158 0.0325158
R3688 AVDD.n683 AVDD.n663 0.0320529
R3689 AVDD.n685 AVDD.n684 0.0320529
R3690 AVDD.n1098 AVDD.n1097 0.0320529
R3691 AVDD.n942 AVDD.n941 0.0320529
R3692 AVDD.n945 AVDD.n944 0.0320529
R3693 AVDD.n943 AVDD.n918 0.0320529
R3694 AVDD.n1027 AVDD.n1026 0.0320529
R3695 AVDD.n1377 AVDD.n1371 0.0319413
R3696 AVDD.n1377 AVDD.n1376 0.0319104
R3697 AVDD.n1122 AVDD.n1121 0.0319052
R3698 AVDD.n1120 AVDD.n1119 0.0319052
R3699 AVDD.n693 AVDD.n665 0.0319052
R3700 AVDD.n1155 AVDD.n56 0.031686
R3701 AVDD.n1157 AVDD.n1156 0.031686
R3702 AVDD.n1159 AVDD.n1158 0.031686
R3703 AVDD.n1216 AVDD.n1215 0.031686
R3704 AVDD.n1214 AVDD.n1213 0.031686
R3705 AVDD.n746 AVDD.n745 0.031686
R3706 AVDD.n744 AVDD.n659 0.031686
R3707 AVDD.n1152 AVDD.n1151 0.031686
R3708 AVDD.n1150 AVDD.n1149 0.031686
R3709 AVDD.n1148 AVDD.n1147 0.031686
R3710 AVDD.n1211 AVDD.n1210 0.031686
R3711 AVDD.n1209 AVDD.n1208 0.031686
R3712 AVDD.n1206 AVDD.n1205 0.031686
R3713 AVDD.n1204 AVDD.n653 0.031686
R3714 AVDD.n1225 AVDD.n1224 0.031686
R3715 AVDD.n1223 AVDD.n1222 0.031686
R3716 AVDD.n747 AVDD.n654 0.031686
R3717 AVDD.n749 AVDD.n748 0.031686
R3718 AVDD.n387 AVDD.n386 0.0315742
R3719 AVDD.n379 AVDD.n378 0.0315742
R3720 AVDD.n536 AVDD.n535 0.0315742
R3721 AVDD.n528 AVDD.n527 0.0315742
R3722 AVDD.n1983 AVDD.n1982 0.0315742
R3723 AVDD.n854 AVDD.n853 0.0315742
R3724 AVDD.n1355 AVDD.n1354 0.0315707
R3725 AVDD.n1360 AVDD.n1359 0.0315707
R3726 AVDD.n1370 AVDD.n1369 0.0315707
R3727 AVDD.n1375 AVDD.n1374 0.0315707
R3728 AVDD.n2010 AVDD.n2009 0.0315707
R3729 AVDD.n2005 AVDD.n2004 0.0315707
R3730 AVDD.n1996 AVDD.n1995 0.0315707
R3731 AVDD.n1407 AVDD.n1401 0.0313793
R3732 AVDD.n1412 AVDD.n1411 0.0313793
R3733 AVDD.n442 AVDD.n440 0.0313793
R3734 AVDD.n510 AVDD.n508 0.0313793
R3735 AVDD.n826 AVDD.n824 0.0313793
R3736 AVDD.n840 AVDD.n839 0.0313793
R3737 AVDD.n1949 AVDD.n1942 0.0313793
R3738 AVDD.n1954 AVDD.n1953 0.0313793
R3739 AVDD.n1143 AVDD.n1142 0.0311937
R3740 AVDD.n311 AVDD.n310 0.0309082
R3741 AVDD.n313 AVDD.n312 0.0309082
R3742 AVDD.n315 AVDD.n314 0.0309082
R3743 AVDD.n319 AVDD.n318 0.0309082
R3744 AVDD.n321 AVDD.n320 0.0309082
R3745 AVDD.n346 AVDD.n345 0.0309082
R3746 AVDD.n348 AVDD.n347 0.0309082
R3747 AVDD.n352 AVDD.n351 0.0309082
R3748 AVDD.n354 AVDD.n353 0.0309082
R3749 AVDD.n561 AVDD.n560 0.0309082
R3750 AVDD.n559 AVDD.n558 0.0309082
R3751 AVDD.n463 AVDD.n462 0.0309082
R3752 AVDD.n465 AVDD.n464 0.0309082
R3753 AVDD.n468 AVDD.n467 0.0309082
R3754 AVDD.n466 AVDD.n356 0.0309082
R3755 AVDD.n551 AVDD.n550 0.0309082
R3756 AVDD.n549 AVDD.n548 0.0309082
R3757 AVDD.n547 AVDD.n546 0.0309082
R3758 AVDD.n1768 AVDD.n1767 0.0303814
R3759 AVDD.n1437 AVDD.n82 0.0303814
R3760 AVDD.n1623 AVDD.n1622 0.0303814
R3761 AVDD.n164 AVDD.n163 0.0303814
R3762 AVDD.n1783 AVDD.n1782 0.0302628
R3763 AVDD.n1452 AVDD.n1451 0.0302628
R3764 AVDD.n1935 AVDD.n43 0.0302628
R3765 AVDD.n1604 AVDD.n66 0.0302628
R3766 AVDD.n1011 AVDD.n1010 0.0295514
R3767 AVDD.n384 AVDD.n383 0.0295026
R3768 AVDD.n533 AVDD.n532 0.0295026
R3769 AVDD.n1980 AVDD.n1979 0.0295026
R3770 AVDD.n553 AVDD.n552 0.0293776
R3771 AVDD.n976 AVDD.n975 0.0289485
R3772 AVDD.n316 AVDD.n315 0.0273367
R3773 AVDD.n988 AVDD.n930 0.0261926
R3774 AVDD.n933 AVDD.n932 0.0259774
R3775 AVDD.n973 AVDD.n972 0.0234742
R3776 AVDD.n975 AVDD.n974 0.0234742
R3777 AVDD.n1418 AVDD.n102 0.0228966
R3778 AVDD.n502 AVDD.n448 0.0228966
R3779 AVDD.n833 AVDD.n832 0.0228966
R3780 AVDD.n1960 AVDD.n33 0.0228966
R3781 AVDD.n1418 AVDD.n1417 0.0228448
R3782 AVDD.n503 AVDD.n502 0.0228448
R3783 AVDD.n834 AVDD.n833 0.0228448
R3784 AVDD.n1960 AVDD.n1959 0.0228448
R3785 AVDD.n985 AVDD.n984 0.0224615
R3786 AVDD.n2018 AVDD.n2 0.0217183
R3787 AVDD.n1366 AVDD.n1365 0.0217183
R3788 AVDD.n2014 AVDD.n2013 0.0217183
R3789 AVDD.n2000 AVDD.n1999 0.0217183
R3790 AVDD.n1400 AVDD.n1399 0.0206724
R3791 AVDD.n1405 AVDD.n1404 0.0206724
R3792 AVDD.n1414 AVDD.n1413 0.0206724
R3793 AVDD.n123 AVDD.n122 0.0206724
R3794 AVDD.n439 AVDD.n438 0.0206724
R3795 AVDD.n445 AVDD.n444 0.0206724
R3796 AVDD.n507 AVDD.n506 0.0206724
R3797 AVDD.n513 AVDD.n512 0.0206724
R3798 AVDD.n823 AVDD.n822 0.0206724
R3799 AVDD.n829 AVDD.n828 0.0206724
R3800 AVDD.n838 AVDD.n837 0.0206724
R3801 AVDD.n843 AVDD.n842 0.0206724
R3802 AVDD.n1941 AVDD.n1940 0.0206724
R3803 AVDD.n1947 AVDD.n1946 0.0206724
R3804 AVDD.n1956 AVDD.n1955 0.0206724
R3805 AVDD.n1260 AVDD.n1259 0.0206724
R3806 AVDD.n1780 AVDD.n54 0.0204161
R3807 AVDD.n1449 AVDD.n77 0.0204161
R3808 AVDD.n1933 AVDD.n1932 0.0204161
R3809 AVDD.n1602 AVDD.n1601 0.0204161
R3810 AVDD.n1756 AVDD.n62 0.019782
R3811 AVDD.n295 AVDD.n142 0.019782
R3812 AVDD.n1634 AVDD.n64 0.019782
R3813 AVDD.n175 AVDD.n146 0.019782
R3814 AVDD.n342 AVDD.n341 0.0196477
R3815 AVDD.n472 AVDD.n471 0.0196477
R3816 AVDD.n753 AVDD.n752 0.0196477
R3817 AVDD.n1202 AVDD.n1201 0.0196477
R3818 AVDD.n2019 AVDD.n2018 0.0189386
R3819 AVDD.n1365 AVDD.n1363 0.0189386
R3820 AVDD.n2014 AVDD.n10 0.0189386
R3821 AVDD.n2001 AVDD.n2000 0.0189386
R3822 AVDD.n959 AVDD.n958 0.0185
R3823 AVDD AVDD.n2022 0.0182591
R3824 AVDD.n991 AVDD.n930 0.0179831
R3825 AVDD.n967 AVDD.n933 0.0178367
R3826 AVDD.n1757 AVDD.n1756 0.0177463
R3827 AVDD.n307 AVDD.n295 0.0177463
R3828 AVDD.n1634 AVDD.n1633 0.0177463
R3829 AVDD.n175 AVDD.n174 0.0177463
R3830 AVDD.n1357 AVDD.n1311 0.0174226
R3831 AVDD.n1961 AVDD.n1960 0.0174226
R3832 AVDD.n502 AVDD.n437 0.0174226
R3833 AVDD.n2007 AVDD.n12 0.0174226
R3834 AVDD.n1418 AVDD.n101 0.0174226
R3835 AVDD.n1357 AVDD.n1351 0.0174226
R3836 AVDD.n1419 AVDD.n1418 0.0174226
R3837 AVDD.n502 AVDD.n501 0.0174226
R3838 AVDD.n833 AVDD.n780 0.0174226
R3839 AVDD.n2007 AVDD.n13 0.0174226
R3840 AVDD.n833 AVDD.n821 0.0174226
R3841 AVDD.n1960 AVDD.n32 0.0174226
R3842 AVDD.n1311 AVDD.n1293 0.0171298
R3843 AVDD.n1309 AVDD.n1293 0.0171298
R3844 AVDD.n1309 AVDD.n1308 0.0171298
R3845 AVDD.n1308 AVDD.n1307 0.0171298
R3846 AVDD.n1307 AVDD.n1296 0.0171298
R3847 AVDD.n1304 AVDD.n1296 0.0171298
R3848 AVDD.n1304 AVDD.n1303 0.0171298
R3849 AVDD.n1303 AVDD.n1302 0.0171298
R3850 AVDD.n1301 AVDD.n1299 0.0171298
R3851 AVDD.n1299 AVDD.n24 0.0171298
R3852 AVDD.n1974 AVDD.n1973 0.0171298
R3853 AVDD.n1973 AVDD.n26 0.0171298
R3854 AVDD.n1971 AVDD.n26 0.0171298
R3855 AVDD.n1970 AVDD.n27 0.0171298
R3856 AVDD.n1968 AVDD.n27 0.0171298
R3857 AVDD.n1968 AVDD.n1967 0.0171298
R3858 AVDD.n1967 AVDD.n1966 0.0171298
R3859 AVDD.n1966 AVDD.n30 0.0171298
R3860 AVDD.n1963 AVDD.n30 0.0171298
R3861 AVDD.n1963 AVDD.n1962 0.0171298
R3862 AVDD.n1962 AVDD.n1961 0.0171298
R3863 AVDD.n437 AVDD.n397 0.0171298
R3864 AVDD.n435 AVDD.n397 0.0171298
R3865 AVDD.n435 AVDD.n434 0.0171298
R3866 AVDD.n434 AVDD.n433 0.0171298
R3867 AVDD.n433 AVDD.n400 0.0171298
R3868 AVDD.n430 AVDD.n400 0.0171298
R3869 AVDD.n430 AVDD.n429 0.0171298
R3870 AVDD.n429 AVDD.n428 0.0171298
R3871 AVDD.n427 AVDD.n402 0.0171298
R3872 AVDD.n425 AVDD.n402 0.0171298
R3873 AVDD.n423 AVDD.n422 0.0171298
R3874 AVDD.n422 AVDD.n405 0.0171298
R3875 AVDD.n420 AVDD.n405 0.0171298
R3876 AVDD.n419 AVDD.n406 0.0171298
R3877 AVDD.n417 AVDD.n406 0.0171298
R3878 AVDD.n417 AVDD.n416 0.0171298
R3879 AVDD.n416 AVDD.n415 0.0171298
R3880 AVDD.n415 AVDD.n409 0.0171298
R3881 AVDD.n412 AVDD.n409 0.0171298
R3882 AVDD.n412 AVDD.n411 0.0171298
R3883 AVDD.n411 AVDD.n12 0.0171298
R3884 AVDD.n1322 AVDD.n101 0.0171298
R3885 AVDD.n1324 AVDD.n1322 0.0171298
R3886 AVDD.n1324 AVDD.n1321 0.0171298
R3887 AVDD.n1327 AVDD.n1321 0.0171298
R3888 AVDD.n1327 AVDD.n1320 0.0171298
R3889 AVDD.n1330 AVDD.n1320 0.0171298
R3890 AVDD.n1330 AVDD.n1319 0.0171298
R3891 AVDD.n1332 AVDD.n1319 0.0171298
R3892 AVDD.n1333 AVDD.n1318 0.0171298
R3893 AVDD.n1335 AVDD.n1318 0.0171298
R3894 AVDD.n1338 AVDD.n1317 0.0171298
R3895 AVDD.n1338 AVDD.n1316 0.0171298
R3896 AVDD.n1340 AVDD.n1316 0.0171298
R3897 AVDD.n1341 AVDD.n1315 0.0171298
R3898 AVDD.n1343 AVDD.n1315 0.0171298
R3899 AVDD.n1343 AVDD.n1314 0.0171298
R3900 AVDD.n1346 AVDD.n1314 0.0171298
R3901 AVDD.n1346 AVDD.n1313 0.0171298
R3902 AVDD.n1349 AVDD.n1313 0.0171298
R3903 AVDD.n1349 AVDD.n1312 0.0171298
R3904 AVDD.n1351 AVDD.n1312 0.0171298
R3905 AVDD.n343 AVDD.n342 0.0171298
R3906 AVDD.n341 AVDD.n323 0.0171298
R3907 AVDD.n339 AVDD.n323 0.0171298
R3908 AVDD.n339 AVDD.n338 0.0171298
R3909 AVDD.n338 AVDD.n337 0.0171298
R3910 AVDD.n337 AVDD.n326 0.0171298
R3911 AVDD.n334 AVDD.n326 0.0171298
R3912 AVDD.n334 AVDD.n333 0.0171298
R3913 AVDD.n333 AVDD.n332 0.0171298
R3914 AVDD.n331 AVDD.n329 0.0171298
R3915 AVDD.n329 AVDD.n93 0.0171298
R3916 AVDD.n1432 AVDD.n1431 0.0171298
R3917 AVDD.n1431 AVDD.n95 0.0171298
R3918 AVDD.n1429 AVDD.n95 0.0171298
R3919 AVDD.n1428 AVDD.n96 0.0171298
R3920 AVDD.n1426 AVDD.n96 0.0171298
R3921 AVDD.n1426 AVDD.n1425 0.0171298
R3922 AVDD.n1425 AVDD.n1424 0.0171298
R3923 AVDD.n1424 AVDD.n99 0.0171298
R3924 AVDD.n1421 AVDD.n99 0.0171298
R3925 AVDD.n1421 AVDD.n1420 0.0171298
R3926 AVDD.n1420 AVDD.n1419 0.0171298
R3927 AVDD.n471 AVDD.n461 0.0171298
R3928 AVDD.n472 AVDD.n460 0.0171298
R3929 AVDD.n474 AVDD.n460 0.0171298
R3930 AVDD.n474 AVDD.n459 0.0171298
R3931 AVDD.n477 AVDD.n459 0.0171298
R3932 AVDD.n477 AVDD.n458 0.0171298
R3933 AVDD.n480 AVDD.n458 0.0171298
R3934 AVDD.n480 AVDD.n457 0.0171298
R3935 AVDD.n482 AVDD.n457 0.0171298
R3936 AVDD.n483 AVDD.n455 0.0171298
R3937 AVDD.n485 AVDD.n455 0.0171298
R3938 AVDD.n488 AVDD.n454 0.0171298
R3939 AVDD.n488 AVDD.n453 0.0171298
R3940 AVDD.n490 AVDD.n453 0.0171298
R3941 AVDD.n491 AVDD.n452 0.0171298
R3942 AVDD.n493 AVDD.n452 0.0171298
R3943 AVDD.n493 AVDD.n451 0.0171298
R3944 AVDD.n496 AVDD.n451 0.0171298
R3945 AVDD.n496 AVDD.n450 0.0171298
R3946 AVDD.n499 AVDD.n450 0.0171298
R3947 AVDD.n499 AVDD.n449 0.0171298
R3948 AVDD.n501 AVDD.n449 0.0171298
R3949 AVDD.n780 AVDD.n729 0.0171298
R3950 AVDD.n778 AVDD.n729 0.0171298
R3951 AVDD.n778 AVDD.n777 0.0171298
R3952 AVDD.n777 AVDD.n776 0.0171298
R3953 AVDD.n776 AVDD.n732 0.0171298
R3954 AVDD.n773 AVDD.n732 0.0171298
R3955 AVDD.n773 AVDD.n772 0.0171298
R3956 AVDD.n772 AVDD.n771 0.0171298
R3957 AVDD.n770 AVDD.n734 0.0171298
R3958 AVDD.n768 AVDD.n734 0.0171298
R3959 AVDD.n766 AVDD.n765 0.0171298
R3960 AVDD.n765 AVDD.n737 0.0171298
R3961 AVDD.n763 AVDD.n737 0.0171298
R3962 AVDD.n762 AVDD.n738 0.0171298
R3963 AVDD.n760 AVDD.n738 0.0171298
R3964 AVDD.n760 AVDD.n759 0.0171298
R3965 AVDD.n759 AVDD.n758 0.0171298
R3966 AVDD.n758 AVDD.n741 0.0171298
R3967 AVDD.n755 AVDD.n741 0.0171298
R3968 AVDD.n755 AVDD.n754 0.0171298
R3969 AVDD.n754 AVDD.n753 0.0171298
R3970 AVDD.n752 AVDD.n743 0.0171298
R3971 AVDD.n792 AVDD.n13 0.0171298
R3972 AVDD.n794 AVDD.n792 0.0171298
R3973 AVDD.n794 AVDD.n791 0.0171298
R3974 AVDD.n797 AVDD.n791 0.0171298
R3975 AVDD.n797 AVDD.n790 0.0171298
R3976 AVDD.n800 AVDD.n790 0.0171298
R3977 AVDD.n800 AVDD.n789 0.0171298
R3978 AVDD.n802 AVDD.n789 0.0171298
R3979 AVDD.n803 AVDD.n787 0.0171298
R3980 AVDD.n805 AVDD.n787 0.0171298
R3981 AVDD.n808 AVDD.n786 0.0171298
R3982 AVDD.n808 AVDD.n785 0.0171298
R3983 AVDD.n810 AVDD.n785 0.0171298
R3984 AVDD.n811 AVDD.n784 0.0171298
R3985 AVDD.n813 AVDD.n784 0.0171298
R3986 AVDD.n813 AVDD.n783 0.0171298
R3987 AVDD.n816 AVDD.n783 0.0171298
R3988 AVDD.n816 AVDD.n782 0.0171298
R3989 AVDD.n819 AVDD.n782 0.0171298
R3990 AVDD.n819 AVDD.n781 0.0171298
R3991 AVDD.n821 AVDD.n781 0.0171298
R3992 AVDD.n1172 AVDD.n32 0.0171298
R3993 AVDD.n1174 AVDD.n1172 0.0171298
R3994 AVDD.n1174 AVDD.n1171 0.0171298
R3995 AVDD.n1177 AVDD.n1171 0.0171298
R3996 AVDD.n1177 AVDD.n1170 0.0171298
R3997 AVDD.n1180 AVDD.n1170 0.0171298
R3998 AVDD.n1180 AVDD.n1169 0.0171298
R3999 AVDD.n1182 AVDD.n1169 0.0171298
R4000 AVDD.n1183 AVDD.n1167 0.0171298
R4001 AVDD.n1185 AVDD.n1167 0.0171298
R4002 AVDD.n1188 AVDD.n1166 0.0171298
R4003 AVDD.n1188 AVDD.n1165 0.0171298
R4004 AVDD.n1190 AVDD.n1165 0.0171298
R4005 AVDD.n1191 AVDD.n1164 0.0171298
R4006 AVDD.n1193 AVDD.n1164 0.0171298
R4007 AVDD.n1193 AVDD.n1163 0.0171298
R4008 AVDD.n1196 AVDD.n1163 0.0171298
R4009 AVDD.n1196 AVDD.n1162 0.0171298
R4010 AVDD.n1199 AVDD.n1162 0.0171298
R4011 AVDD.n1199 AVDD.n1161 0.0171298
R4012 AVDD.n1201 AVDD.n1161 0.0171298
R4013 AVDD.n1202 AVDD.n1160 0.0171298
R4014 AVDD.n322 AVDD.n141 0.0166614
R4015 AVDD.n470 AVDD.n357 0.0166614
R4016 AVDD.n981 AVDD.n980 0.0163144
R4017 AVDD.n1302 AVDD.n1301 0.01631
R4018 AVDD.n1971 AVDD.n1970 0.01631
R4019 AVDD.n428 AVDD.n427 0.01631
R4020 AVDD.n420 AVDD.n419 0.01631
R4021 AVDD.n1333 AVDD.n1332 0.01631
R4022 AVDD.n1341 AVDD.n1340 0.01631
R4023 AVDD.n332 AVDD.n331 0.01631
R4024 AVDD.n1429 AVDD.n1428 0.01631
R4025 AVDD.n483 AVDD.n482 0.01631
R4026 AVDD.n491 AVDD.n490 0.01631
R4027 AVDD.n771 AVDD.n770 0.01631
R4028 AVDD.n763 AVDD.n762 0.01631
R4029 AVDD.n803 AVDD.n802 0.01631
R4030 AVDD.n811 AVDD.n810 0.01631
R4031 AVDD.n1183 AVDD.n1182 0.01631
R4032 AVDD.n1191 AVDD.n1190 0.01631
R4033 AVDD.n55 AVDD.n54 0.0162238
R4034 AVDD.n78 AVDD.n77 0.0162238
R4035 AVDD.n1932 AVDD.n45 0.0162238
R4036 AVDD.n1601 AVDD.n68 0.0162238
R4037 AVDD.n1397 AVDD.n1396 0.0159138
R4038 AVDD.n1399 AVDD.n1398 0.0159138
R4039 AVDD.n1401 AVDD.n1400 0.0159138
R4040 AVDD.n1406 AVDD.n1405 0.0159138
R4041 AVDD.n1404 AVDD.n1403 0.0159138
R4042 AVDD.n1402 AVDD.n102 0.0159138
R4043 AVDD.n1417 AVDD.n1416 0.0159138
R4044 AVDD.n1415 AVDD.n1414 0.0159138
R4045 AVDD.n1413 AVDD.n1412 0.0159138
R4046 AVDD.n122 AVDD.n103 0.0159138
R4047 AVDD.n124 AVDD.n123 0.0159138
R4048 AVDD.n438 AVDD.n125 0.0159138
R4049 AVDD.n440 AVDD.n439 0.0159138
R4050 AVDD.n444 AVDD.n443 0.0159138
R4051 AVDD.n446 AVDD.n445 0.0159138
R4052 AVDD.n448 AVDD.n447 0.0159138
R4053 AVDD.n504 AVDD.n503 0.0159138
R4054 AVDD.n506 AVDD.n505 0.0159138
R4055 AVDD.n508 AVDD.n507 0.0159138
R4056 AVDD.n512 AVDD.n511 0.0159138
R4057 AVDD.n514 AVDD.n513 0.0159138
R4058 AVDD.n516 AVDD.n515 0.0159138
R4059 AVDD.n822 AVDD.n635 0.0159138
R4060 AVDD.n824 AVDD.n823 0.0159138
R4061 AVDD.n828 AVDD.n827 0.0159138
R4062 AVDD.n830 AVDD.n829 0.0159138
R4063 AVDD.n832 AVDD.n831 0.0159138
R4064 AVDD.n835 AVDD.n834 0.0159138
R4065 AVDD.n837 AVDD.n836 0.0159138
R4066 AVDD.n839 AVDD.n838 0.0159138
R4067 AVDD.n842 AVDD.n841 0.0159138
R4068 AVDD.n844 AVDD.n843 0.0159138
R4069 AVDD.n1938 AVDD.n1937 0.0159138
R4070 AVDD.n1940 AVDD.n1939 0.0159138
R4071 AVDD.n1942 AVDD.n1941 0.0159138
R4072 AVDD.n1948 AVDD.n1947 0.0159138
R4073 AVDD.n1946 AVDD.n1945 0.0159138
R4074 AVDD.n1944 AVDD.n33 0.0159138
R4075 AVDD.n1959 AVDD.n1958 0.0159138
R4076 AVDD.n1957 AVDD.n1956 0.0159138
R4077 AVDD.n1955 AVDD.n1954 0.0159138
R4078 AVDD.n1259 AVDD.n34 0.0159138
R4079 AVDD.n1261 AVDD.n1260 0.0159138
R4080 AVDD.n983 AVDD.n982 0.0156839
R4081 AVDD.n980 AVDD.n977 0.0154737
R4082 AVDD.n1975 AVDD.n24 0.015256
R4083 AVDD.n425 AVDD.n424 0.015256
R4084 AVDD.n1335 AVDD.n110 0.015256
R4085 AVDD.n1433 AVDD.n93 0.015256
R4086 AVDD.n485 AVDD.n456 0.015256
R4087 AVDD.n768 AVDD.n767 0.015256
R4088 AVDD.n805 AVDD.n788 0.015256
R4089 AVDD.n1185 AVDD.n1168 0.015256
R4090 AVDD.n1051 AVDD.n1050 0.0148793
R4091 AVDD.n935 AVDD.n899 0.0142069
R4092 AVDD.n1357 AVDD.n1356 0.0138734
R4093 AVDD.n2008 AVDD.n2007 0.0138734
R4094 AVDD.n926 AVDD.n925 0.0138448
R4095 AVDD.n1358 AVDD.n1357 0.0138425
R4096 AVDD.n2007 AVDD.n2006 0.0138425
R4097 AVDD AVDD.n0 0.0138116
R4098 AVDD.n860 AVDD.n859 0.012725
R4099 AVDD.n2021 AVDD.n2020 0.0125453
R4100 AVDD.n1353 AVDD.n1352 0.0125453
R4101 AVDD.n1362 AVDD.n1361 0.0125453
R4102 AVDD.n1368 AVDD.n1367 0.0125453
R4103 AVDD.n1373 AVDD.n1372 0.0125453
R4104 AVDD.n2012 AVDD.n2011 0.0125453
R4105 AVDD.n2003 AVDD.n2002 0.0125453
R4106 AVDD.n1998 AVDD.n1997 0.0125453
R4107 AVDD.n977 AVDD.n976 0.0119536
R4108 AVDD.n982 AVDD.n981 0.0119536
R4109 AVDD.n984 AVDD.n983 0.0119536
R4110 AVDD.n961 AVDD.n960 0.0117759
R4111 AVDD.n940 AVDD.n939 0.0117759
R4112 AVDD.n1049 AVDD.n1048 0.0117759
R4113 AVDD.n925 AVDD.n900 0.0117759
R4114 AVDD.n987 AVDD.n986 0.0116909
R4115 AVDD.n565 AVDD.n564 0.0113718
R4116 AVDD.n595 AVDD.n594 0.0113718
R4117 AVDD.n600 AVDD.n599 0.0113718
R4118 AVDD.n1265 AVDD.n1264 0.0113718
R4119 AVDD.n1257 AVDD.n1256 0.0113718
R4120 AVDD.n1229 AVDD.n1228 0.0113718
R4121 AVDD.n938 AVDD.n937 0.0111034
R4122 AVDD.n751 AVDD.n750 0.0108058
R4123 AVDD.n1212 AVDD.n1203 0.0108058
R4124 AVDD.n344 AVDD.n322 0.0101617
R4125 AVDD.n470 AVDD.n469 0.0101617
R4126 AVDD.n1378 AVDD.n1377 0.0101084
R4127 AVDD.n1377 AVDD.n1292 0.0101084
R4128 AVDD.n564 AVDD.n139 0.00994219
R4129 AVDD.n565 AVDD.n138 0.00994219
R4130 AVDD.n567 AVDD.n138 0.00994219
R4131 AVDD.n567 AVDD.n137 0.00994219
R4132 AVDD.n570 AVDD.n137 0.00994219
R4133 AVDD.n570 AVDD.n136 0.00994219
R4134 AVDD.n573 AVDD.n136 0.00994219
R4135 AVDD.n573 AVDD.n135 0.00994219
R4136 AVDD.n575 AVDD.n135 0.00994219
R4137 AVDD.n576 AVDD.n133 0.00994219
R4138 AVDD.n578 AVDD.n133 0.00994219
R4139 AVDD.n581 AVDD.n132 0.00994219
R4140 AVDD.n581 AVDD.n131 0.00994219
R4141 AVDD.n583 AVDD.n131 0.00994219
R4142 AVDD.n584 AVDD.n130 0.00994219
R4143 AVDD.n586 AVDD.n130 0.00994219
R4144 AVDD.n586 AVDD.n129 0.00994219
R4145 AVDD.n589 AVDD.n129 0.00994219
R4146 AVDD.n589 AVDD.n128 0.00994219
R4147 AVDD.n592 AVDD.n128 0.00994219
R4148 AVDD.n592 AVDD.n127 0.00994219
R4149 AVDD.n594 AVDD.n127 0.00994219
R4150 AVDD.n595 AVDD.n126 0.00994219
R4151 AVDD.n596 AVDD.n126 0.00994219
R4152 AVDD.n598 AVDD.n121 0.00994219
R4153 AVDD.n599 AVDD.n121 0.00994219
R4154 AVDD.n600 AVDD.n120 0.00994219
R4155 AVDD.n602 AVDD.n120 0.00994219
R4156 AVDD.n602 AVDD.n119 0.00994219
R4157 AVDD.n605 AVDD.n119 0.00994219
R4158 AVDD.n605 AVDD.n118 0.00994219
R4159 AVDD.n608 AVDD.n118 0.00994219
R4160 AVDD.n608 AVDD.n117 0.00994219
R4161 AVDD.n610 AVDD.n117 0.00994219
R4162 AVDD.n613 AVDD.n612 0.00994219
R4163 AVDD.n612 AVDD.n114 0.00994219
R4164 AVDD.n1391 AVDD.n1390 0.00994219
R4165 AVDD.n1390 AVDD.n116 0.00994219
R4166 AVDD.n1388 AVDD.n116 0.00994219
R4167 AVDD.n1387 AVDD.n615 0.00994219
R4168 AVDD.n1385 AVDD.n615 0.00994219
R4169 AVDD.n1385 AVDD.n1384 0.00994219
R4170 AVDD.n1384 AVDD.n1383 0.00994219
R4171 AVDD.n1383 AVDD.n618 0.00994219
R4172 AVDD.n1380 AVDD.n618 0.00994219
R4173 AVDD.n1380 AVDD.n1379 0.00994219
R4174 AVDD.n1379 AVDD.n1378 0.00994219
R4175 AVDD.n1292 AVDD.n620 0.00994219
R4176 AVDD.n1290 AVDD.n620 0.00994219
R4177 AVDD.n1290 AVDD.n1289 0.00994219
R4178 AVDD.n1289 AVDD.n1288 0.00994219
R4179 AVDD.n1288 AVDD.n623 0.00994219
R4180 AVDD.n1285 AVDD.n623 0.00994219
R4181 AVDD.n1285 AVDD.n1284 0.00994219
R4182 AVDD.n1284 AVDD.n1283 0.00994219
R4183 AVDD.n1282 AVDD.n625 0.00994219
R4184 AVDD.n1280 AVDD.n625 0.00994219
R4185 AVDD.n1278 AVDD.n1277 0.00994219
R4186 AVDD.n1277 AVDD.n628 0.00994219
R4187 AVDD.n1275 AVDD.n628 0.00994219
R4188 AVDD.n1274 AVDD.n629 0.00994219
R4189 AVDD.n1272 AVDD.n629 0.00994219
R4190 AVDD.n1272 AVDD.n1271 0.00994219
R4191 AVDD.n1271 AVDD.n1270 0.00994219
R4192 AVDD.n1270 AVDD.n632 0.00994219
R4193 AVDD.n1267 AVDD.n632 0.00994219
R4194 AVDD.n1267 AVDD.n1266 0.00994219
R4195 AVDD.n1266 AVDD.n1265 0.00994219
R4196 AVDD.n1264 AVDD.n634 0.00994219
R4197 AVDD.n1263 AVDD.n634 0.00994219
R4198 AVDD.n1258 AVDD.n636 0.00994219
R4199 AVDD.n1257 AVDD.n636 0.00994219
R4200 AVDD.n1256 AVDD.n637 0.00994219
R4201 AVDD.n1254 AVDD.n637 0.00994219
R4202 AVDD.n1254 AVDD.n1253 0.00994219
R4203 AVDD.n1253 AVDD.n1252 0.00994219
R4204 AVDD.n1252 AVDD.n640 0.00994219
R4205 AVDD.n1249 AVDD.n640 0.00994219
R4206 AVDD.n1249 AVDD.n1248 0.00994219
R4207 AVDD.n1248 AVDD.n1247 0.00994219
R4208 AVDD.n1246 AVDD.n642 0.00994219
R4209 AVDD.n1244 AVDD.n642 0.00994219
R4210 AVDD.n1242 AVDD.n1241 0.00994219
R4211 AVDD.n1241 AVDD.n646 0.00994219
R4212 AVDD.n1239 AVDD.n646 0.00994219
R4213 AVDD.n1238 AVDD.n647 0.00994219
R4214 AVDD.n1236 AVDD.n647 0.00994219
R4215 AVDD.n1236 AVDD.n1235 0.00994219
R4216 AVDD.n1235 AVDD.n1234 0.00994219
R4217 AVDD.n1234 AVDD.n650 0.00994219
R4218 AVDD.n1231 AVDD.n650 0.00994219
R4219 AVDD.n1231 AVDD.n1230 0.00994219
R4220 AVDD.n1230 AVDD.n1229 0.00994219
R4221 AVDD.n1228 AVDD.n652 0.00994219
R4222 AVDD.n1605 AVDD.n0 0.00970384
R4223 AVDD.n2022 AVDD.n2021 0.00970384
R4224 AVDD.n2020 AVDD.n2019 0.00970384
R4225 AVDD.n1352 AVDD.n2 0.00970384
R4226 AVDD.n1354 AVDD.n1353 0.00970384
R4227 AVDD.n1356 AVDD.n1355 0.00970384
R4228 AVDD.n1359 AVDD.n1358 0.00970384
R4229 AVDD.n1361 AVDD.n1360 0.00970384
R4230 AVDD.n1363 AVDD.n1362 0.00970384
R4231 AVDD.n1367 AVDD.n1366 0.00970384
R4232 AVDD.n1369 AVDD.n1368 0.00970384
R4233 AVDD.n1371 AVDD.n1370 0.00970384
R4234 AVDD.n1376 AVDD.n1375 0.00970384
R4235 AVDD.n1374 AVDD.n1373 0.00970384
R4236 AVDD.n1372 AVDD.n10 0.00970384
R4237 AVDD.n2013 AVDD.n2012 0.00970384
R4238 AVDD.n2011 AVDD.n2010 0.00970384
R4239 AVDD.n2009 AVDD.n2008 0.00970384
R4240 AVDD.n2006 AVDD.n2005 0.00970384
R4241 AVDD.n2004 AVDD.n2003 0.00970384
R4242 AVDD.n2002 AVDD.n2001 0.00970384
R4243 AVDD.n1999 AVDD.n1998 0.00970384
R4244 AVDD.n1997 AVDD.n1996 0.00970384
R4245 AVDD.n1995 AVDD.n1994 0.00970384
R4246 AVDD.n563 AVDD.n140 0.00967621
R4247 AVDD.n576 AVDD.n575 0.00947673
R4248 AVDD.n584 AVDD.n583 0.00947673
R4249 AVDD.n613 AVDD.n610 0.00947673
R4250 AVDD.n1388 AVDD.n1387 0.00947673
R4251 AVDD.n1283 AVDD.n1282 0.00947673
R4252 AVDD.n1275 AVDD.n1274 0.00947673
R4253 AVDD.n1247 AVDD.n1246 0.00947673
R4254 AVDD.n1239 AVDD.n1238 0.00947673
R4255 AVDD.n1047 AVDD.n900 0.00944828
R4256 AVDD.n597 AVDD.n596 0.00927724
R4257 AVDD.n598 AVDD.n597 0.00927724
R4258 AVDD.n1263 AVDD.n1262 0.00927724
R4259 AVDD.n1262 AVDD.n1258 0.00927724
R4260 AVDD.n578 AVDD.n134 0.00887828
R4261 AVDD.n1392 AVDD.n114 0.00887828
R4262 AVDD.n1280 AVDD.n1279 0.00887828
R4263 AVDD.n1244 AVDD.n1243 0.00887828
R4264 AVDD.n927 AVDD.n926 0.00877586
R4265 AVDD.n1096 AVDD.n686 0.00791176
R4266 AVDD.n1061 AVDD.n1060 0.00787705
R4267 AVDD.n928 AVDD.n927 0.00763793
R4268 AVDD.n344 AVDD.n343 0.00746812
R4269 AVDD.n469 AVDD.n461 0.00746812
R4270 AVDD.n884 AVDD.n883 0.0073513
R4271 AVDD.n726 AVDD.n725 0.0073513
R4272 AVDD.n697 AVDD.n696 0.0073513
R4273 AVDD.n890 AVDD.n698 0.0073513
R4274 AVDD.n889 AVDD.n888 0.0073513
R4275 AVDD.n702 AVDD.n700 0.0073513
R4276 AVDD.n721 AVDD.n720 0.0073513
R4277 AVDD.n717 AVDD.n706 0.0073513
R4278 AVDD.n716 AVDD.n715 0.0073513
R4279 AVDD.n714 AVDD.n707 0.0073513
R4280 AVDD.n887 AVDD.n723 0.00713029
R4281 AVDD.n703 AVDD.n699 0.00713029
R4282 AVDD.n881 AVDD.n727 0.0070075
R4283 AVDD.n880 AVDD.n724 0.0070075
R4284 AVDD.n710 AVDD.n709 0.0070075
R4285 AVDD.n712 AVDD.n711 0.0070075
R4286 AVDD.n936 AVDD.n935 0.00696552
R4287 AVDD.n863 AVDD.n862 0.00693383
R4288 AVDD.n866 AVDD.n848 0.00693383
R4289 AVDD.n869 AVDD.n867 0.00693383
R4290 AVDD.n868 AVDD.n846 0.00693383
R4291 AVDD.n871 AVDD.n870 0.00693383
R4292 AVDD.n750 AVDD.n743 0.00682401
R4293 AVDD.n1212 AVDD.n1160 0.00682401
R4294 AVDD.n704 AVDD.n701 0.00656548
R4295 AVDD.n894 AVDD.n695 0.00651637
R4296 AVDD.n1048 AVDD.n1047 0.0065
R4297 AVDD.n847 AVDD.n845 0.0064427
R4298 AVDD.n1227 AVDD.n1226 0.0063515
R4299 AVDD.n563 AVDD.n562 0.00598578
R4300 AVDD.n876 AVDD.n874 0.00595157
R4301 AVDD.n875 AVDD.n728 0.00595157
R4302 AVDD.n878 AVDD.n877 0.00595157
R4303 AVDD.n1139 AVDD.n662 0.00595157
R4304 AVDD.n1142 AVDD.n661 0.00595157
R4305 AVDD.n937 AVDD.n936 0.00531034
R4306 AVDD.n1012 AVDD.n1011 0.00512451
R4307 AVDD.n350 AVDD.n349 0.00509184
R4308 AVDD.n557 AVDD.n355 0.00509184
R4309 AVDD.n858 AVDD.n664 0.00489563
R4310 AVDD.n939 AVDD.n938 0.00484483
R4311 AVDD.n562 AVDD.n139 0.00445641
R4312 AVDD.n1783 AVDD.n55 0.00441304
R4313 AVDD.n1452 AVDD.n78 0.00441304
R4314 AVDD.n45 AVDD.n43 0.00441304
R4315 AVDD.n68 AVDD.n66 0.00441304
R4316 AVDD.n1769 AVDD.n1768 0.00429447
R4317 AVDD.n1438 AVDD.n1437 0.00429447
R4318 AVDD.n1622 AVDD.n1621 0.00429447
R4319 AVDD.n163 AVDD.n162 0.00429447
R4320 AVDD.n383 AVDD.n382 0.00418286
R4321 AVDD.n532 AVDD.n531 0.00418286
R4322 AVDD.n1979 AVDD.n19 0.00418286
R4323 AVDD.n1226 AVDD.n652 0.00409069
R4324 AVDD.n958 AVDD.n940 0.00355172
R4325 AVDD.n1137 AVDD.n1136 0.00342224
R4326 AVDD.n517 AVDD.n516 0.00334483
R4327 AVDD.n1138 AVDD.n1137 0.00302933
R4328 AVDD.n997 AVDD.n928 0.00277586
R4329 AVDD.n1396 AVDD.n79 0.00272414
R4330 AVDD.n1937 AVDD.n1936 0.00272414
R4331 AVDD.n962 AVDD.n961 0.00267241
R4332 AVDD.n864 AVDD.n664 0.0025382
R4333 AVDD.n1975 AVDD.n1974 0.00237378
R4334 AVDD.n424 AVDD.n423 0.00237378
R4335 AVDD.n1317 AVDD.n110 0.00237378
R4336 AVDD.n1433 AVDD.n1432 0.00237378
R4337 AVDD.n456 AVDD.n454 0.00237378
R4338 AVDD.n767 AVDD.n766 0.00237378
R4339 AVDD.n788 AVDD.n786 0.00237378
R4340 AVDD.n1168 AVDD.n1166 0.00237378
R4341 AVDD.n997 AVDD.n996 0.00236207
R4342 AVDD.n1994 AVDD.n1993 0.0021987
R4343 AVDD.n867 AVDD.n866 0.00209618
R4344 AVDD.n876 AVDD.n875 0.00202251
R4345 AVDD.n878 AVDD.n728 0.00202251
R4346 AVDD.n877 AVDD.n727 0.00202251
R4347 AVDD.n711 AVDD.n662 0.00202251
R4348 AVDD.n1139 AVDD.n1138 0.00202251
R4349 AVDD.n1136 AVDD.n661 0.00202251
R4350 AVDD.n962 AVDD.n694 0.00189655
R4351 AVDD.n1606 AVDD.n1605 0.00182807
R4352 AVDD.n1050 AVDD.n1049 0.00168966
R4353 AVDD.n1904 AVDD.n1903 0.00168421
R4354 AVDD.n1899 AVDD.n1898 0.00168421
R4355 AVDD.n1894 AVDD.n1893 0.00168421
R4356 AVDD.n1889 AVDD.n1888 0.00168421
R4357 AVDD.n1807 AVDD.n1806 0.00168421
R4358 AVDD.n1802 AVDD.n1801 0.00168421
R4359 AVDD.n1797 AVDD.n1796 0.00168421
R4360 AVDD.n1856 AVDD.n1855 0.00168421
R4361 AVDD.n1851 AVDD.n1850 0.00168421
R4362 AVDD.n1846 AVDD.n1845 0.00168421
R4363 AVDD.n1841 AVDD.n1840 0.00168421
R4364 AVDD.n1826 AVDD.n1825 0.00168421
R4365 AVDD.n1821 AVDD.n1820 0.00168421
R4366 AVDD.n1816 AVDD.n1815 0.00168421
R4367 AVDD.n1651 AVDD.n1648 0.00168421
R4368 AVDD.n1660 AVDD.n1658 0.00168421
R4369 AVDD.n1663 AVDD.n1655 0.00168421
R4370 AVDD.n1645 AVDD.n1642 0.00168421
R4371 AVDD.n1709 AVDD.n1640 0.00168421
R4372 AVDD.n1712 AVDD.n1637 0.00168421
R4373 AVDD.n1563 AVDD.n1485 0.00168421
R4374 AVDD.n1566 AVDD.n1482 0.00168421
R4375 AVDD.n1569 AVDD.n1479 0.00168421
R4376 AVDD.n1572 AVDD.n1476 0.00168421
R4377 AVDD.n1472 AVDD.n1471 0.00168421
R4378 AVDD.n1467 AVDD.n1466 0.00168421
R4379 AVDD.n1462 AVDD.n1461 0.00168421
R4380 AVDD.n1523 AVDD.n1522 0.00168421
R4381 AVDD.n1526 AVDD.n1519 0.00168421
R4382 AVDD.n1529 AVDD.n1516 0.00168421
R4383 AVDD.n1532 AVDD.n1513 0.00168421
R4384 AVDD.n1509 AVDD.n1508 0.00168421
R4385 AVDD.n1504 AVDD.n1503 0.00168421
R4386 AVDD.n1499 AVDD.n1498 0.00168421
R4387 AVDD.n209 AVDD.n206 0.00168421
R4388 AVDD.n203 AVDD.n202 0.00168421
R4389 AVDD.n198 AVDD.n197 0.00168421
R4390 AVDD.n252 AVDD.n249 0.00168421
R4391 AVDD.n246 AVDD.n245 0.00168421
R4392 AVDD.n241 AVDD.n240 0.00168421
R4393 AVDD.n1101 AVDD.n682 0.00168421
R4394 AVDD.n1104 AVDD.n679 0.00168421
R4395 AVDD.n1107 AVDD.n676 0.00168421
R4396 AVDD.n1110 AVDD.n673 0.00168421
R4397 AVDD.n1113 AVDD.n671 0.00168421
R4398 AVDD.n1116 AVDD.n668 0.00168421
R4399 AVDD.n1094 AVDD.n1092 0.00168421
R4400 AVDD.n1088 AVDD.n1086 0.00168421
R4401 AVDD.n1082 AVDD.n1080 0.00168421
R4402 AVDD.n1076 AVDD.n1075 0.00168421
R4403 AVDD.n1072 AVDD.n1070 0.00168421
R4404 AVDD.n1066 AVDD.n1064 0.00168421
R4405 AVDD.n1030 AVDD.n917 0.00168421
R4406 AVDD.n1033 AVDD.n914 0.00168421
R4407 AVDD.n1036 AVDD.n911 0.00168421
R4408 AVDD.n1039 AVDD.n908 0.00168421
R4409 AVDD.n1042 AVDD.n906 0.00168421
R4410 AVDD.n1045 AVDD.n903 0.00168421
R4411 AVDD.n134 AVDD.n132 0.00156391
R4412 AVDD.n1392 AVDD.n1391 0.00156391
R4413 AVDD.n1279 AVDD.n1278 0.00156391
R4414 AVDD.n1243 AVDD.n1242 0.00156391
R4415 AVDD.n1051 AVDD.n899 0.00153448
R4416 AVDD.n874 AVDD.n845 0.00153138
R4417 AVDD.n894 AVDD.n893 0.00133493
R4418 AVDD.n705 AVDD.n704 0.00128581
R4419 AVDD.n960 AVDD.n959 0.00106897
R4420 AVDD.n859 AVDD.n858 0.00104025
R4421 AVDD.n864 AVDD.n863 0.00104025
R4422 AVDD.n862 AVDD.n848 0.00104025
R4423 AVDD.n869 AVDD.n868 0.00104025
R4424 AVDD.n871 AVDD.n846 0.00104025
R4425 AVDD.n870 AVDD.n847 0.00104025
R4426 AVDD.n881 AVDD.n880 0.000966576
R4427 AVDD.n712 AVDD.n710 0.000966576
R4428 AVDD.n987 AVDD.n985 0.000762697
R4429 AVDD.n723 AVDD.n699 0.00072101
R4430 AVDD.n884 AVDD.n724 0.000622783
R4431 AVDD.n883 AVDD.n726 0.000622783
R4432 AVDD.n725 AVDD.n695 0.000622783
R4433 AVDD.n893 AVDD.n696 0.000622783
R4434 AVDD.n698 AVDD.n697 0.000622783
R4435 AVDD.n890 AVDD.n889 0.000622783
R4436 AVDD.n888 AVDD.n887 0.000622783
R4437 AVDD.n703 AVDD.n702 0.000622783
R4438 AVDD.n721 AVDD.n700 0.000622783
R4439 AVDD.n720 AVDD.n701 0.000622783
R4440 AVDD.n706 AVDD.n705 0.000622783
R4441 AVDD.n717 AVDD.n716 0.000622783
R4442 AVDD.n715 AVDD.n714 0.000622783
R4443 AVDD.n709 AVDD.n707 0.000622783
R4444 AVSS.n172 AVSS.n171 4252.69
R4445 AVSS.n438 AVSS.n437 661.869
R4446 AVSS.n394 AVSS.n175 661.869
R4447 AVSS.n391 AVSS.n62 661.869
R4448 AVSS.n64 AVSS.n63 656.895
R4449 AVSS.n434 AVSS.n173 656.895
R4450 AVSS.n441 AVSS.n61 656.895
R4451 AVSS.n437 AVSS.n64 656.434
R4452 AVSS.n434 AVSS.n175 656.434
R4453 AVSS.n441 AVSS.n62 656.434
R4454 AVSS.n438 AVSS.n63 653.672
R4455 AVSS.n394 AVSS.n173 653.672
R4456 AVSS.n391 AVSS.n61 653.672
R4457 AVSS.t31 AVSS.t79 517.433
R4458 AVSS.t46 AVSS.t138 517.433
R4459 AVSS.t98 AVSS.t1 454.447
R4460 AVSS.t28 AVSS.t178 450.327
R4461 AVSS.n107 AVSS.n78 383.618
R4462 AVSS.n147 AVSS.n78 381.962
R4463 AVSS.n107 AVSS.n77 381.132
R4464 AVSS.n147 AVSS.n77 379.474
R4465 AVSS.t133 AVSS.t31 329.651
R4466 AVSS.t138 AVSS.t95 329.651
R4467 AVSS.n107 AVSS.t46 275.635
R4468 AVSS.n171 AVSS.t1 275.495
R4469 AVSS.n149 AVSS.t28 275.495
R4470 AVSS.n148 AVSS.t79 275.495
R4471 AVSS.n150 AVSS.n67 267.474
R4472 AVSS.n170 AVSS.n67 266.829
R4473 AVSS.n150 AVSS.n66 266.276
R4474 AVSS.n170 AVSS.n66 265.632
R4475 AVSS.t95 AVSS.n106 244.294
R4476 AVSS.n106 AVSS.t133 233.7
R4477 AVSS.t235 AVSS.t74 178.191
R4478 AVSS.t172 AVSS.t43 178.191
R4479 AVSS.t144 AVSS.t201 173.123
R4480 AVSS.t16 AVSS.t175 173.123
R4481 AVSS.t178 AVSS.n76 168.946
R4482 AVSS.n76 AVSS.t98 160.706
R4483 AVSS.t55 AVSS.t158 158.528
R4484 AVSS.t64 AVSS.t25 158.528
R4485 AVSS.t85 AVSS.t114 155.487
R4486 AVSS.t10 AVSS.t22 155.487
R4487 AVSS.t7 AVSS.t235 113.523
R4488 AVSS.t201 AVSS.t7 113.523
R4489 AVSS.t222 AVSS.t144 113.523
R4490 AVSS.t175 AVSS.t40 113.523
R4491 AVSS.t40 AVSS.t172 113.523
R4492 AVSS.n435 AVSS.t16 109.469
R4493 AVSS.t13 AVSS.t163 95.8869
R4494 AVSS.t103 AVSS.t82 95.8869
R4495 AVSS.t74 AVSS.n391 94.9497
R4496 AVSS.t43 AVSS.n172 94.8732
R4497 AVSS.t67 AVSS.t19 93.8597
R4498 AVSS.t4 AVSS.t155 93.8597
R4499 AVSS.t34 AVSS.t52 90.8189
R4500 AVSS.n174 AVSS.t49 89.6025
R4501 AVSS.n149 AVSS.n148 84.7678
R4502 AVSS.n393 AVSS.t141 80.2775
R4503 AVSS.n440 AVSS.t88 80.2775
R4504 AVSS.n393 AVSS.n392 32.0302
R4505 AVSS.n440 AVSS.n439 29.1921
R4506 AVSS.t49 AVSS.t85 22.7051
R4507 AVSS.t22 AVSS.t34 22.7051
R4508 AVSS.t158 AVSS.t67 19.6643
R4509 AVSS.t19 AVSS.t4 19.6643
R4510 AVSS.t155 AVSS.t64 19.6643
R4511 AVSS.t114 AVSS.t13 17.6371
R4512 AVSS.t163 AVSS.t103 17.6371
R4513 AVSS.t82 AVSS.t10 17.6371
R4514 AVSS.t141 AVSS.t55 14.5963
R4515 AVSS.t25 AVSS.t88 14.5963
R4516 AVSS.n156 AVSS.t118 8.52542
R4517 AVSS.n79 AVSS.t78 8.52542
R4518 AVSS.n111 AVSS.t182 8.52542
R4519 AVSS.n115 AVSS.t213 8.52542
R4520 AVSS.n90 AVSS.t137 8.52542
R4521 AVSS.n98 AVSS.t94 8.52542
R4522 AVSS.n91 AVSS.t132 8.52542
R4523 AVSS.n92 AVSS.t211 8.52542
R4524 AVSS.n103 AVSS.t245 8.52542
R4525 AVSS.n105 AVSS.t203 8.52542
R4526 AVSS.n137 AVSS.t45 8.52542
R4527 AVSS.n135 AVSS.t71 8.52542
R4528 AVSS.n109 AVSS.t247 8.52542
R4529 AVSS.n130 AVSS.t180 8.52542
R4530 AVSS.n110 AVSS.t241 8.52542
R4531 AVSS.n124 AVSS.t30 8.52542
R4532 AVSS.n491 AVSS.t148 8.06917
R4533 AVSS.n222 AVSS.t9 8.06917
R4534 AVSS.n214 AVSS.t102 8.06917
R4535 AVSS.n212 AVSS.t12 8.06917
R4536 AVSS.n233 AVSS.t84 8.06917
R4537 AVSS.n207 AVSS.t165 8.06917
R4538 AVSS.n201 AVSS.t87 8.06917
R4539 AVSS.n244 AVSS.t63 8.06917
R4540 AVSS.n197 AVSS.t146 8.06917
R4541 AVSS.n195 AVSS.t66 8.06917
R4542 AVSS.n192 AVSS.t251 8.06917
R4543 AVSS.n2 AVSS.t51 8.06917
R4544 AVSS.n216 AVSS.t263 8.06917
R4545 AVSS.n223 AVSS.t81 8.06917
R4546 AVSS.n213 AVSS.t162 8.06917
R4547 AVSS.n211 AVSS.t113 8.06917
R4548 AVSS.n234 AVSS.t167 8.06917
R4549 AVSS.n200 AVSS.t76 8.06917
R4550 AVSS.n245 AVSS.t154 8.06917
R4551 AVSS.n196 AVSS.t259 8.06917
R4552 AVSS.n194 AVSS.t157 8.06917
R4553 AVSS.n191 AVSS.t140 8.06917
R4554 AVSS.n204 AVSS.t48 8.06917
R4555 AVSS.n203 AVSS.t111 8.06917
R4556 AVSS.n444 AVSS.t275 8.06917
R4557 AVSS.n445 AVSS.t126 8.06917
R4558 AVSS.n447 AVSS.t215 8.06917
R4559 AVSS.n204 AVSS.t230 8.06917
R4560 AVSS.n203 AVSS.t271 8.06917
R4561 AVSS.n444 AVSS.t184 8.06917
R4562 AVSS.n445 AVSS.t24 8.06917
R4563 AVSS.n447 AVSS.t116 8.06917
R4564 AVSS.n280 AVSS.t205 8.06917
R4565 AVSS.n284 AVSS.t18 8.06917
R4566 AVSS.n279 AVSS.t207 8.06917
R4567 AVSS.n278 AVSS.t188 8.06917
R4568 AVSS.n292 AVSS.t257 8.06917
R4569 AVSS.n277 AVSS.t190 8.06917
R4570 AVSS.n276 AVSS.t243 8.06917
R4571 AVSS.n299 AVSS.t69 8.06917
R4572 AVSS.n275 AVSS.t267 8.06917
R4573 AVSS.n351 AVSS.t224 8.06917
R4574 AVSS.n354 AVSS.t39 8.06917
R4575 AVSS.n350 AVSS.t226 8.06917
R4576 AVSS.n359 AVSS.t15 8.06917
R4577 AVSS.n362 AVSS.t105 8.06917
R4578 AVSS.n349 AVSS.t21 8.06917
R4579 AVSS.n348 AVSS.t120 8.06917
R4580 AVSS.n369 AVSS.t209 8.06917
R4581 AVSS.n347 AVSS.t130 8.06917
R4582 AVSS.n9 AVSS.t124 8.06917
R4583 AVSS.n475 AVSS.t92 8.06917
R4584 AVSS.n5 AVSS.t171 8.06917
R4585 AVSS.n480 AVSS.t269 8.06917
R4586 AVSS.n4 AVSS.t174 8.06917
R4587 AVSS.n485 AVSS.t261 8.06917
R4588 AVSS.n6 AVSS.t237 8.06917
R4589 AVSS.n6 AVSS.t281 8.06917
R4590 AVSS.n6 AVSS.t194 8.06917
R4591 AVSS.n6 AVSS.t42 8.06917
R4592 AVSS.n400 AVSS.t122 8.06917
R4593 AVSS.n398 AVSS.t273 8.06917
R4594 AVSS.n397 AVSS.t135 8.06917
R4595 AVSS.n187 AVSS.t54 8.06917
R4596 AVSS.n188 AVSS.t160 8.06917
R4597 AVSS.n176 AVSS.t150 8.06917
R4598 AVSS.n420 AVSS.t232 8.06917
R4599 AVSS.n177 AVSS.t152 8.06917
R4600 AVSS.n178 AVSS.t217 8.06917
R4601 AVSS.n412 AVSS.t36 8.06917
R4602 AVSS.n179 AVSS.t219 8.06917
R4603 AVSS.n180 AVSS.t196 8.06917
R4604 AVSS.n405 AVSS.t3 8.06917
R4605 AVSS.n181 AVSS.t198 8.06917
R4606 AVSS.n425 AVSS.t33 8.06917
R4607 AVSS.n427 AVSS.t192 8.06917
R4608 AVSS.n428 AVSS.t59 8.06917
R4609 AVSS.n431 AVSS.t239 8.06917
R4610 AVSS.n430 AVSS.t90 8.06917
R4611 AVSS.n258 AVSS.t221 8.06917
R4612 AVSS.n185 AVSS.t143 8.06917
R4613 AVSS.n184 AVSS.t200 8.06917
R4614 AVSS.n265 AVSS.t6 8.06917
R4615 AVSS.n183 AVSS.t234 8.06917
R4616 AVSS.n270 AVSS.t128 8.06917
R4617 AVSS.n272 AVSS.t279 8.06917
R4618 AVSS.n273 AVSS.t73 8.06917
R4619 AVSS.n388 AVSS.t249 8.06917
R4620 AVSS.n387 AVSS.t107 8.06917
R4621 AVSS.n385 AVSS.t169 8.06917
R4622 AVSS.n319 AVSS.t313 6.72766
R4623 AVSS.n69 AVSS.t0 6.60917
R4624 AVSS.n69 AVSS.t253 6.60917
R4625 AVSS.n69 AVSS.t61 6.60917
R4626 AVSS.n69 AVSS.t100 6.60917
R4627 AVSS.n69 AVSS.t277 6.60917
R4628 AVSS.n162 AVSS.t186 6.60917
R4629 AVSS.n72 AVSS.t109 6.60917
R4630 AVSS.n116 AVSS.t177 6.60917
R4631 AVSS.n71 AVSS.t97 6.60917
R4632 AVSS.n157 AVSS.t265 6.60917
R4633 AVSS.n154 AVSS.t228 6.60917
R4634 AVSS.n75 AVSS.t27 6.60917
R4635 AVSS.n80 AVSS.t57 6.60917
R4636 AVSS.n112 AVSS.t255 6.60917
R4637 AVSS.n34 AVSS.t344 6.53862
R4638 AVSS.n70 AVSS.t333 5.49372
R4639 AVSS.n317 AVSS.t342 5.47432
R4640 AVSS.n312 AVSS.n311 5.31981
R4641 AVSS.n38 AVSS.t306 5.28484
R4642 AVSS.n43 AVSS.t302 5.28484
R4643 AVSS.n37 AVSS.t285 5.28484
R4644 AVSS.n316 AVSS.n303 5.26136
R4645 AVSS.t2 AVSS.n167 5.2505
R4646 AVSS.n168 AVSS.t2 5.2505
R4647 AVSS.n167 AVSS.t254 5.2505
R4648 AVSS.n168 AVSS.t254 5.2505
R4649 AVSS.n167 AVSS.t62 5.2505
R4650 AVSS.n168 AVSS.t62 5.2505
R4651 AVSS.n167 AVSS.t101 5.2505
R4652 AVSS.n168 AVSS.t101 5.2505
R4653 AVSS.n167 AVSS.t278 5.2505
R4654 AVSS.n168 AVSS.t278 5.2505
R4655 AVSS.n161 AVSS.t187 5.2505
R4656 AVSS.n165 AVSS.t110 5.2505
R4657 AVSS.t99 AVSS.n70 5.2505
R4658 AVSS.n120 AVSS.t179 5.2505
R4659 AVSS.n56 AVSS.n55 5.16888
R4660 AVSS.n20 AVSS.n19 5.15456
R4661 AVSS.n376 AVSS.n375 5.09675
R4662 AVSS.n464 AVSS.n461 4.63106
R4663 AVSS.n455 AVSS.n452 4.63106
R4664 AVSS.n27 AVSS.n24 4.63106
R4665 AVSS.n313 AVSS.n312 4.61712
R4666 AVSS.n380 AVSS.n379 4.61712
R4667 AVSS.n141 AVSS.n140 4.61585
R4668 AVSS.n144 AVSS.n143 4.61585
R4669 AVSS.n378 AVSS.n377 4.61078
R4670 AVSS.n468 AVSS.n466 4.61078
R4671 AVSS.n459 AVSS.n457 4.61078
R4672 AVSS.n31 AVSS.n29 4.61078
R4673 AVSS.n22 AVSS.n20 4.61078
R4674 AVSS.n377 AVSS.n376 4.60825
R4675 AVSS.n469 AVSS.n468 4.60825
R4676 AVSS.n460 AVSS.n459 4.60825
R4677 AVSS.n32 AVSS.n31 4.60825
R4678 AVSS.n23 AVSS.n22 4.60825
R4679 AVSS.n320 AVSS.n317 4.60439
R4680 AVSS.n140 AVSS.n139 4.60318
R4681 AVSS.n143 AVSS.n142 4.60318
R4682 AVSS.n314 AVSS.n313 4.60191
R4683 AVSS.n381 AVSS.n380 4.60191
R4684 AVSS.n465 AVSS.n464 4.58796
R4685 AVSS.n456 AVSS.n455 4.58796
R4686 AVSS.n28 AVSS.n27 4.58796
R4687 AVSS.n305 AVSS.n304 4.5005
R4688 AVSS.n308 AVSS.n306 4.5005
R4689 AVSS.n310 AVSS.n309 4.5005
R4690 AVSS.n21 AVSS.n18 4.5005
R4691 AVSS.n26 AVSS.n17 4.5005
R4692 AVSS.n30 AVSS.n16 4.5005
R4693 AVSS.n454 AVSS.n15 4.5005
R4694 AVSS.n458 AVSS.n14 4.5005
R4695 AVSS.n463 AVSS.n13 4.5005
R4696 AVSS.n467 AVSS.n12 4.5005
R4697 AVSS.n84 AVSS.n82 4.5005
R4698 AVSS.n88 AVSS.n86 4.5005
R4699 AVSS.n333 AVSS.t327 4.41563
R4700 AVSS.n342 AVSS.t340 4.41563
R4701 AVSS.n331 AVSS.t311 4.41563
R4702 AVSS.n321 AVSS.t360 4.41563
R4703 AVSS.n50 AVSS.t295 4.22616
R4704 AVSS.n48 AVSS.t354 4.22616
R4705 AVSS.n319 AVSS.n318 4.21432
R4706 AVSS.n316 AVSS.n315 4.21432
R4707 AVSS.n439 AVSS.t37 4.05489
R4708 AVSS.n40 AVSS.n39 4.02484
R4709 AVSS.n42 AVSS.n41 4.02484
R4710 AVSS.n36 AVSS.n35 4.02484
R4711 AVSS.n34 AVSS.n33 4.02484
R4712 AVSS.n50 AVSS.t288 4.02247
R4713 AVSS.n48 AVSS.t300 4.02247
R4714 AVSS.n310 AVSS.t349 4.00471
R4715 AVSS.n305 AVSS.t346 4.00471
R4716 AVSS.n51 AVSS.n11 3.96014
R4717 AVSS.n333 AVSS.t304 3.833
R4718 AVSS.n342 AVSS.t348 3.833
R4719 AVSS.n331 AVSS.t322 3.833
R4720 AVSS.n321 AVSS.t356 3.833
R4721 AVSS.n467 AVSS.t292 3.81405
R4722 AVSS.n458 AVSS.t343 3.81405
R4723 AVSS.n30 AVSS.t325 3.81405
R4724 AVSS.n21 AVSS.t329 3.81405
R4725 AVSS.n330 AVSS.n326 3.80578
R4726 AVSS.n341 AVSS.n337 3.80578
R4727 AVSS.n36 AVSS.n34 3.80578
R4728 AVSS.n42 AVSS.n40 3.80578
R4729 AVSS.n382 AVSS.n381 3.76738
R4730 AVSS.n473 AVSS.t125 3.37683
R4731 AVSS.t149 AVSS.n1 3.3605
R4732 AVSS.n217 AVSS.t149 3.3605
R4733 AVSS.n219 AVSS.t11 3.3605
R4734 AVSS.t14 AVSS.n210 3.3605
R4735 AVSS.n231 AVSS.t86 3.3605
R4736 AVSS.t89 AVSS.n199 3.3605
R4737 AVSS.n241 AVSS.t65 3.3605
R4738 AVSS.t68 AVSS.n193 3.3605
R4739 AVSS.n253 AVSS.t252 3.3605
R4740 AVSS.t252 AVSS.n186 3.3605
R4741 AVSS.n218 AVSS.t264 3.3605
R4742 AVSS.n221 AVSS.t83 3.3605
R4743 AVSS.n230 AVSS.t115 3.3605
R4744 AVSS.n232 AVSS.t168 3.3605
R4745 AVSS.t168 AVSS.n209 3.3605
R4746 AVSS.t77 AVSS.n239 3.3605
R4747 AVSS.n240 AVSS.t77 3.3605
R4748 AVSS.n243 AVSS.t156 3.3605
R4749 AVSS.n252 AVSS.t159 3.3605
R4750 AVSS.t142 AVSS.n254 3.3605
R4751 AVSS.t206 AVSS.n281 3.3605
R4752 AVSS.n287 AVSS.t208 3.3605
R4753 AVSS.t189 AVSS.n288 3.3605
R4754 AVSS.n295 AVSS.t191 3.3605
R4755 AVSS.t244 AVSS.n296 3.3605
R4756 AVSS.n302 AVSS.t268 3.3605
R4757 AVSS.t225 AVSS.n10 3.3605
R4758 AVSS.n357 AVSS.t227 3.3605
R4759 AVSS.n358 AVSS.t17 3.3605
R4760 AVSS.n365 AVSS.t23 3.3605
R4761 AVSS.t121 AVSS.n366 3.3605
R4762 AVSS.n372 AVSS.t131 3.3605
R4763 AVSS.t125 AVSS.n472 3.3605
R4764 AVSS.t173 AVSS.n477 3.3605
R4765 AVSS.n483 AVSS.t176 3.3605
R4766 AVSS.n484 AVSS.t262 3.3605
R4767 AVSS.n8 AVSS.t282 3.3605
R4768 AVSS.t282 AVSS.n7 3.3605
R4769 AVSS.n8 AVSS.t195 3.3605
R4770 AVSS.n7 AVSS.t195 3.3605
R4771 AVSS.n8 AVSS.t44 3.3605
R4772 AVSS.n7 AVSS.t44 3.3605
R4773 AVSS.n423 AVSS.t151 3.3605
R4774 AVSS.t153 AVSS.n417 3.3605
R4775 AVSS.n416 AVSS.t218 3.3605
R4776 AVSS.t220 AVSS.n409 3.3605
R4777 AVSS.n408 AVSS.t197 3.3605
R4778 AVSS.t199 AVSS.n402 3.3605
R4779 AVSS.n261 AVSS.t145 3.3605
R4780 AVSS.t202 AVSS.n262 3.3605
R4781 AVSS.n268 AVSS.t236 3.3605
R4782 AVSS.n336 AVSS.n334 3.15563
R4783 AVSS.n340 AVSS.n338 3.15563
R4784 AVSS.n329 AVSS.n327 3.15563
R4785 AVSS.n325 AVSS.n323 3.15563
R4786 AVSS.n119 AVSS.n118 3.1505
R4787 AVSS.n164 AVSS.n163 3.1505
R4788 AVSS.n320 AVSS.n319 3.02463
R4789 AVSS.n54 AVSS.n52 2.96616
R4790 AVSS.n47 AVSS.n45 2.96616
R4791 AVSS.n24 AVSS.n23 2.885
R4792 AVSS.n461 AVSS.n460 2.885
R4793 AVSS.n436 AVSS.n435 2.83857
R4794 AVSS.n452 AVSS.n451 2.795
R4795 AVSS.n54 AVSS.n53 2.76247
R4796 AVSS.n47 AVSS.n46 2.76247
R4797 AVSS.n308 AVSS.n307 2.74471
R4798 AVSS.n49 AVSS.n47 2.71914
R4799 AVSS.n337 AVSS.n333 2.71872
R4800 AVSS.n101 AVSS.t139 2.6955
R4801 AVSS.n97 AVSS.t96 2.6955
R4802 AVSS.n95 AVSS.t134 2.6955
R4803 AVSS.t212 AVSS.n74 2.6955
R4804 AVSS.n133 AVSS.t248 2.6955
R4805 AVSS.n129 AVSS.t181 2.6955
R4806 AVSS.n127 AVSS.t242 2.6955
R4807 AVSS.n123 AVSS.t32 2.6955
R4808 AVSS.n160 AVSS.t266 2.6255
R4809 AVSS.n155 AVSS.t229 2.6255
R4810 AVSS.n153 AVSS.t29 2.6255
R4811 AVSS.n81 AVSS.t58 2.6255
R4812 AVSS.n114 AVSS.t256 2.6255
R4813 AVSS.n336 AVSS.n335 2.573
R4814 AVSS.n340 AVSS.n339 2.573
R4815 AVSS.n329 AVSS.n328 2.573
R4816 AVSS.n325 AVSS.n324 2.573
R4817 AVSS.n463 AVSS.n462 2.55405
R4818 AVSS.n454 AVSS.n453 2.55405
R4819 AVSS.n26 AVSS.n25 2.55405
R4820 AVSS.n56 AVSS.n49 2.46014
R4821 AVSS.n145 AVSS.n144 2.45973
R4822 AVSS.n139 AVSS.n138 2.45073
R4823 AVSS.n344 AVSS.n332 2.38034
R4824 AVSS.n38 AVSS.n11 2.37491
R4825 AVSS.n44 AVSS.n43 2.32143
R4826 AVSS.n449 AVSS.n448 2.30076
R4827 AVSS.n375 AVSS.n314 2.26738
R4828 AVSS.n345 AVSS.n320 2.23722
R4829 AVSS.n88 AVSS.n87 2.15932
R4830 AVSS.n84 AVSS.n83 2.15932
R4831 AVSS.n140 AVSS.n89 2.15458
R4832 AVSS.n143 AVSS.n85 2.15458
R4833 AVSS.n57 AVSS.n44 2.13932
R4834 AVSS.n487 AVSS.n486 2.1005
R4835 AVSS.n482 AVSS.n481 2.1005
R4836 AVSS.n479 AVSS.n478 2.1005
R4837 AVSS.t110 AVSS.n164 2.1005
R4838 AVSS.n164 AVSS.t187 2.1005
R4839 AVSS.n119 AVSS.t99 2.1005
R4840 AVSS.t179 AVSS.n119 2.1005
R4841 AVSS.n404 AVSS.n403 2.1005
R4842 AVSS.n407 AVSS.n406 2.1005
R4843 AVSS.n411 AVSS.n410 2.1005
R4844 AVSS.n415 AVSS.n414 2.1005
R4845 AVSS.n419 AVSS.n418 2.1005
R4846 AVSS.n422 AVSS.n421 2.1005
R4847 AVSS.n267 AVSS.n266 2.1005
R4848 AVSS.n264 AVSS.n263 2.1005
R4849 AVSS.n260 AVSS.n259 2.1005
R4850 AVSS.n371 AVSS.n370 2.1005
R4851 AVSS.n368 AVSS.n367 2.1005
R4852 AVSS.n364 AVSS.n363 2.1005
R4853 AVSS.n361 AVSS.n360 2.1005
R4854 AVSS.n356 AVSS.n355 2.1005
R4855 AVSS.n353 AVSS.n352 2.1005
R4856 AVSS.n301 AVSS.n300 2.1005
R4857 AVSS.n298 AVSS.n297 2.1005
R4858 AVSS.n294 AVSS.n293 2.1005
R4859 AVSS.n290 AVSS.n289 2.1005
R4860 AVSS.n286 AVSS.n285 2.1005
R4861 AVSS.n283 AVSS.n282 2.1005
R4862 AVSS.n256 AVSS.n255 2.1005
R4863 AVSS.n251 AVSS.n250 2.1005
R4864 AVSS.n242 AVSS.n198 2.1005
R4865 AVSS.n229 AVSS.n228 2.1005
R4866 AVSS.n220 AVSS.n215 2.1005
R4867 AVSS.n489 AVSS.n488 2.1005
R4868 AVSS.n249 AVSS.n248 2.1005
R4869 AVSS.n247 AVSS.n246 2.1005
R4870 AVSS.n238 AVSS.n237 2.1005
R4871 AVSS.n236 AVSS.n235 2.1005
R4872 AVSS.n227 AVSS.n226 2.1005
R4873 AVSS.n225 AVSS.n224 2.1005
R4874 AVSS.n471 AVSS.n470 1.7274
R4875 AVSS.n205 AVSS.t50 1.6805
R4876 AVSS.n202 AVSS.t112 1.6805
R4877 AVSS.n443 AVSS.t276 1.6805
R4878 AVSS.n446 AVSS.t127 1.6805
R4879 AVSS.n59 AVSS.t216 1.6805
R4880 AVSS.n205 AVSS.t231 1.6805
R4881 AVSS.n202 AVSS.t272 1.6805
R4882 AVSS.n443 AVSS.t185 1.6805
R4883 AVSS.n446 AVSS.t26 1.6805
R4884 AVSS.n59 AVSS.t117 1.6805
R4885 AVSS.n476 AVSS.t93 1.6805
R4886 AVSS.n474 AVSS.t238 1.6805
R4887 AVSS.n401 AVSS.t123 1.6805
R4888 AVSS.n399 AVSS.t274 1.6805
R4889 AVSS.n396 AVSS.t136 1.6805
R4890 AVSS.n182 AVSS.t56 1.6805
R4891 AVSS.n189 AVSS.t161 1.6805
R4892 AVSS.n424 AVSS.t35 1.6805
R4893 AVSS.n426 AVSS.t193 1.6805
R4894 AVSS.n429 AVSS.t60 1.6805
R4895 AVSS.n432 AVSS.t240 1.6805
R4896 AVSS.n0 AVSS.t91 1.6805
R4897 AVSS.n269 AVSS.t129 1.6805
R4898 AVSS.n271 AVSS.t280 1.6805
R4899 AVSS.n274 AVSS.t75 1.6805
R4900 AVSS.n389 AVSS.t250 1.6805
R4901 AVSS.n386 AVSS.t108 1.6805
R4902 AVSS.n384 AVSS.t170 1.6805
R4903 AVSS.n383 AVSS.n382 1.67828
R4904 AVSS.n374 AVSS.n373 1.67828
R4905 AVSS.n322 AVSS.n303 1.67718
R4906 AVSS.n470 AVSS.n469 1.60175
R4907 AVSS.n126 AVSS.n125 1.5755
R4908 AVSS.n132 AVSS.n131 1.5755
R4909 AVSS.n94 AVSS.n93 1.5755
R4910 AVSS.n100 AVSS.n99 1.5755
R4911 AVSS.n375 AVSS.n374 1.5005
R4912 AVSS.n345 AVSS.n344 1.5005
R4913 AVSS.n451 AVSS.n450 1.5005
R4914 AVSS.n57 AVSS.n56 1.5005
R4915 AVSS.n51 AVSS.n50 1.46537
R4916 AVSS.n55 AVSS.n54 1.46537
R4917 AVSS.n49 AVSS.n48 1.46537
R4918 AVSS.n337 AVSS.n336 1.46537
R4919 AVSS.n341 AVSS.n340 1.46537
R4920 AVSS.n343 AVSS.n342 1.46537
R4921 AVSS.n332 AVSS.n331 1.46537
R4922 AVSS.n330 AVSS.n329 1.46537
R4923 AVSS.n326 AVSS.n325 1.46537
R4924 AVSS.n322 AVSS.n321 1.46537
R4925 AVSS.n158 AVSS.t119 1.348
R4926 AVSS.n152 AVSS.t80 1.348
R4927 AVSS.n113 AVSS.t183 1.348
R4928 AVSS.n122 AVSS.t214 1.348
R4929 AVSS.n102 AVSS.t246 1.348
R4930 AVSS.n104 AVSS.t204 1.348
R4931 AVSS.n136 AVSS.t47 1.348
R4932 AVSS.n134 AVSS.t72 1.348
R4933 AVSS.n142 AVSS.n141 1.265
R4934 AVSS.t104 AVSS.n225 1.2605
R4935 AVSS.n225 AVSS.t11 1.2605
R4936 AVSS.n226 AVSS.t14 1.2605
R4937 AVSS.n226 AVSS.t104 1.2605
R4938 AVSS.t166 AVSS.n236 1.2605
R4939 AVSS.n236 AVSS.t86 1.2605
R4940 AVSS.n237 AVSS.t89 1.2605
R4941 AVSS.n237 AVSS.t166 1.2605
R4942 AVSS.t147 AVSS.n247 1.2605
R4943 AVSS.n247 AVSS.t65 1.2605
R4944 AVSS.n248 AVSS.t68 1.2605
R4945 AVSS.n248 AVSS.t147 1.2605
R4946 AVSS.n488 AVSS.t264 1.2605
R4947 AVSS.n488 AVSS.t53 1.2605
R4948 AVSS.n220 AVSS.t164 1.2605
R4949 AVSS.t83 AVSS.n220 1.2605
R4950 AVSS.t115 AVSS.n229 1.2605
R4951 AVSS.n229 AVSS.t164 1.2605
R4952 AVSS.n242 AVSS.t260 1.2605
R4953 AVSS.t156 AVSS.n242 1.2605
R4954 AVSS.t159 AVSS.n251 1.2605
R4955 AVSS.n251 AVSS.t260 1.2605
R4956 AVSS.n255 AVSS.t223 1.2605
R4957 AVSS.n255 AVSS.t142 1.2605
R4958 AVSS.n282 AVSS.t20 1.2605
R4959 AVSS.n282 AVSS.t206 1.2605
R4960 AVSS.t208 AVSS.n286 1.2605
R4961 AVSS.n286 AVSS.t20 1.2605
R4962 AVSS.n289 AVSS.t258 1.2605
R4963 AVSS.n289 AVSS.t189 1.2605
R4964 AVSS.t191 AVSS.n294 1.2605
R4965 AVSS.n294 AVSS.t258 1.2605
R4966 AVSS.n297 AVSS.t70 1.2605
R4967 AVSS.n297 AVSS.t244 1.2605
R4968 AVSS.t268 AVSS.n301 1.2605
R4969 AVSS.n301 AVSS.t70 1.2605
R4970 AVSS.n352 AVSS.t41 1.2605
R4971 AVSS.n352 AVSS.t225 1.2605
R4972 AVSS.t227 AVSS.n356 1.2605
R4973 AVSS.n356 AVSS.t41 1.2605
R4974 AVSS.t106 AVSS.n361 1.2605
R4975 AVSS.n361 AVSS.t17 1.2605
R4976 AVSS.t23 AVSS.n364 1.2605
R4977 AVSS.n364 AVSS.t106 1.2605
R4978 AVSS.n367 AVSS.t210 1.2605
R4979 AVSS.n367 AVSS.t121 1.2605
R4980 AVSS.t131 AVSS.n371 1.2605
R4981 AVSS.n371 AVSS.t210 1.2605
R4982 AVSS.n311 AVSS.t323 1.2605
R4983 AVSS.n311 AVSS.t351 1.2605
R4984 AVSS.n307 AVSS.t359 1.2605
R4985 AVSS.n307 AVSS.t347 1.2605
R4986 AVSS.n334 AVSS.t326 1.2605
R4987 AVSS.n334 AVSS.t318 1.2605
R4988 AVSS.n335 AVSS.t303 1.2605
R4989 AVSS.n335 AVSS.t328 1.2605
R4990 AVSS.n338 AVSS.t309 1.2605
R4991 AVSS.n338 AVSS.t338 1.2605
R4992 AVSS.n339 AVSS.t339 1.2605
R4993 AVSS.n339 AVSS.t298 1.2605
R4994 AVSS.n327 AVSS.t310 1.2605
R4995 AVSS.n327 AVSS.t296 1.2605
R4996 AVSS.n328 AVSS.t321 1.2605
R4997 AVSS.n328 AVSS.t287 1.2605
R4998 AVSS.n323 AVSS.t335 1.2605
R4999 AVSS.n323 AVSS.t315 1.2605
R5000 AVSS.n324 AVSS.t316 1.2605
R5001 AVSS.n324 AVSS.t286 1.2605
R5002 AVSS.n318 AVSS.t332 1.2605
R5003 AVSS.n318 AVSS.t319 1.2605
R5004 AVSS.n315 AVSS.t341 1.2605
R5005 AVSS.n315 AVSS.t289 1.2605
R5006 AVSS.n52 AVSS.t320 1.2605
R5007 AVSS.n52 AVSS.t301 1.2605
R5008 AVSS.n53 AVSS.t312 1.2605
R5009 AVSS.n53 AVSS.t361 1.2605
R5010 AVSS.n45 AVSS.t290 1.2605
R5011 AVSS.n45 AVSS.t331 1.2605
R5012 AVSS.n46 AVSS.t299 1.2605
R5013 AVSS.n46 AVSS.t307 1.2605
R5014 AVSS.n39 AVSS.t305 1.2605
R5015 AVSS.n39 AVSS.t330 1.2605
R5016 AVSS.n41 AVSS.t283 1.2605
R5017 AVSS.n41 AVSS.t337 1.2605
R5018 AVSS.n35 AVSS.t284 1.2605
R5019 AVSS.n35 AVSS.t314 1.2605
R5020 AVSS.n33 AVSS.t358 1.2605
R5021 AVSS.n33 AVSS.t355 1.2605
R5022 AVSS.n462 AVSS.t291 1.2605
R5023 AVSS.n462 AVSS.t336 1.2605
R5024 AVSS.n453 AVSS.t357 1.2605
R5025 AVSS.n453 AVSS.t293 1.2605
R5026 AVSS.n25 AVSS.t294 1.2605
R5027 AVSS.n25 AVSS.t350 1.2605
R5028 AVSS.n19 AVSS.t297 1.2605
R5029 AVSS.n19 AVSS.t334 1.2605
R5030 AVSS.n478 AVSS.t270 1.2605
R5031 AVSS.n478 AVSS.t173 1.2605
R5032 AVSS.t176 AVSS.n482 1.2605
R5033 AVSS.n482 AVSS.t270 1.2605
R5034 AVSS.t53 AVSS.n487 1.2605
R5035 AVSS.n487 AVSS.t262 1.2605
R5036 AVSS.n422 AVSS.t233 1.2605
R5037 AVSS.t151 AVSS.n422 1.2605
R5038 AVSS.n418 AVSS.t153 1.2605
R5039 AVSS.n418 AVSS.t233 1.2605
R5040 AVSS.n415 AVSS.t38 1.2605
R5041 AVSS.t218 AVSS.n415 1.2605
R5042 AVSS.n410 AVSS.t220 1.2605
R5043 AVSS.n410 AVSS.t38 1.2605
R5044 AVSS.n407 AVSS.t5 1.2605
R5045 AVSS.t197 AVSS.n407 1.2605
R5046 AVSS.n403 AVSS.t199 1.2605
R5047 AVSS.n403 AVSS.t5 1.2605
R5048 AVSS.t145 AVSS.n260 1.2605
R5049 AVSS.n260 AVSS.t223 1.2605
R5050 AVSS.n263 AVSS.t8 1.2605
R5051 AVSS.n263 AVSS.t202 1.2605
R5052 AVSS.t236 AVSS.n267 1.2605
R5053 AVSS.n267 AVSS.t8 1.2605
R5054 AVSS.n326 AVSS.n322 1.25428
R5055 AVSS.n332 AVSS.n330 1.25428
R5056 AVSS.n343 AVSS.n341 1.25428
R5057 AVSS.n317 AVSS.n316 1.25428
R5058 AVSS.n37 AVSS.n36 1.25428
R5059 AVSS.n43 AVSS.n42 1.25428
R5060 AVSS.n40 AVSS.n38 1.25428
R5061 AVSS.n55 AVSS.n51 1.25428
R5062 AVSS.n392 AVSS.t222 1.21682
R5063 AVSS.n174 AVSS.t37 1.21682
R5064 AVSS.n436 AVSS.t52 1.21682
R5065 AVSS.n449 AVSS.n58 1.13691
R5066 AVSS.n100 AVSS.t96 1.1205
R5067 AVSS.t139 AVSS.n100 1.1205
R5068 AVSS.n94 AVSS.t212 1.1205
R5069 AVSS.t134 AVSS.n94 1.1205
R5070 AVSS.n87 AVSS.t308 1.1205
R5071 AVSS.n87 AVSS.t345 1.1205
R5072 AVSS.n89 AVSS.t353 1.1205
R5073 AVSS.n89 AVSS.t363 1.1205
R5074 AVSS.n83 AVSS.t362 1.1205
R5075 AVSS.n83 AVSS.t352 1.1205
R5076 AVSS.n85 AVSS.t324 1.1205
R5077 AVSS.n85 AVSS.t317 1.1205
R5078 AVSS.n132 AVSS.t181 1.1205
R5079 AVSS.t248 AVSS.n132 1.1205
R5080 AVSS.n126 AVSS.t32 1.1205
R5081 AVSS.t242 AVSS.n126 1.1205
R5082 AVSS.n29 AVSS.n28 0.9995
R5083 AVSS.n457 AVSS.n456 0.9995
R5084 AVSS.n466 AVSS.n465 0.9995
R5085 AVSS.n379 AVSS.n378 0.973625
R5086 AVSS.n450 AVSS.n449 0.970331
R5087 AVSS.n382 AVSS.n303 0.585196
R5088 AVSS.n374 AVSS.n345 0.585196
R5089 AVSS.n450 AVSS.n57 0.585196
R5090 AVSS.n470 AVSS.n11 0.585196
R5091 AVSS.n169 AVSS.n68 0.239651
R5092 AVSS.n44 AVSS.n37 0.236091
R5093 AVSS.n151 AVSS.n150 0.186214
R5094 AVSS.n150 AVSS.n149 0.186214
R5095 AVSS.n170 AVSS.n169 0.186214
R5096 AVSS.n171 AVSS.n170 0.186214
R5097 AVSS.n344 AVSS.n343 0.177184
R5098 AVSS.n117 AVSS.n67 0.163
R5099 AVSS.n76 AVSS.n67 0.163
R5100 AVSS.n73 AVSS.n66 0.163
R5101 AVSS.n76 AVSS.n66 0.163
R5102 AVSS.n108 AVSS.n107 0.141041
R5103 AVSS.n147 AVSS.n146 0.141041
R5104 AVSS.n148 AVSS.n147 0.141041
R5105 AVSS.n381 AVSS.n304 0.14
R5106 AVSS.n379 AVSS.n304 0.14
R5107 AVSS.n378 AVSS.n306 0.14
R5108 AVSS.n376 AVSS.n306 0.14
R5109 AVSS.n314 AVSS.n309 0.14
R5110 AVSS.n312 AVSS.n309 0.14
R5111 AVSS.n20 AVSS.n18 0.14
R5112 AVSS.n23 AVSS.n18 0.14
R5113 AVSS.n24 AVSS.n17 0.14
R5114 AVSS.n28 AVSS.n17 0.14
R5115 AVSS.n29 AVSS.n16 0.14
R5116 AVSS.n32 AVSS.n16 0.14
R5117 AVSS.n452 AVSS.n15 0.14
R5118 AVSS.n456 AVSS.n15 0.14
R5119 AVSS.n457 AVSS.n14 0.14
R5120 AVSS.n460 AVSS.n14 0.14
R5121 AVSS.n461 AVSS.n13 0.14
R5122 AVSS.n465 AVSS.n13 0.14
R5123 AVSS.n466 AVSS.n12 0.14
R5124 AVSS.n469 AVSS.n12 0.14
R5125 AVSS.n144 AVSS.n82 0.14
R5126 AVSS.n142 AVSS.n82 0.14
R5127 AVSS.n141 AVSS.n86 0.14
R5128 AVSS.n139 AVSS.n86 0.14
R5129 AVSS.n166 AVSS.n70 0.132207
R5130 AVSS.n128 AVSS.n78 0.108833
R5131 AVSS.n106 AVSS.n78 0.108833
R5132 AVSS.n96 AVSS.n77 0.108833
R5133 AVSS.n106 AVSS.n77 0.108833
R5134 AVSS.n475 AVSS.n474 0.105988
R5135 AVSS.n426 AVSS.n425 0.105988
R5136 AVSS.n400 AVSS.n399 0.105988
R5137 AVSS.n271 AVSS.n270 0.105988
R5138 AVSS.n386 AVSS.n385 0.105988
R5139 AVSS.n490 AVSS.n0 0.102012
R5140 AVSS.n190 AVSS.n189 0.102012
R5141 AVSS.n451 AVSS.n32 0.10175
R5142 AVSS.n166 AVSS.n71 0.100659
R5143 AVSS.n391 AVSS.n390 0.0769706
R5144 AVSS.n395 AVSS.n394 0.0769706
R5145 AVSS.n394 AVSS.n393 0.0769706
R5146 AVSS.n434 AVSS.n433 0.0769706
R5147 AVSS.n435 AVSS.n434 0.0769706
R5148 AVSS.n68 AVSS.n64 0.0769706
R5149 AVSS.n172 AVSS.n64 0.0769706
R5150 AVSS.n442 AVSS.n441 0.0769706
R5151 AVSS.n441 AVSS.n440 0.0769706
R5152 AVSS.n438 AVSS.n60 0.0769706
R5153 AVSS.n439 AVSS.n438 0.0769706
R5154 AVSS.n395 AVSS.n182 0.072814
R5155 AVSS.n390 AVSS.n389 0.072814
R5156 AVSS.n104 AVSS.n103 0.0718609
R5157 AVSS.n136 AVSS.n135 0.0718609
R5158 AVSS.n433 AVSS.n429 0.0681047
R5159 AVSS.n433 AVSS.n432 0.0678953
R5160 AVSS.n257 AVSS.n61 0.0646975
R5161 AVSS.n392 AVSS.n61 0.0646975
R5162 AVSS.n413 AVSS.n173 0.0646975
R5163 AVSS.n174 AVSS.n173 0.0646975
R5164 AVSS.n437 AVSS.n65 0.0646975
R5165 AVSS.n437 AVSS.n436 0.0646975
R5166 AVSS.n291 AVSS.n62 0.0646975
R5167 AVSS.n392 AVSS.n62 0.0646975
R5168 AVSS.n63 AVSS.n3 0.0646975
R5169 AVSS.n436 AVSS.n63 0.0646975
R5170 AVSS.n208 AVSS.n175 0.0646975
R5171 AVSS.n175 AVSS.n174 0.0646975
R5172 AVSS.n396 AVSS.n395 0.063186
R5173 AVSS.n390 AVSS.n274 0.063186
R5174 AVSS.n447 AVSS.n446 0.0533671
R5175 AVSS.n206 AVSS.n205 0.0513741
R5176 AVSS.n165 AVSS.n72 0.0431396
R5177 AVSS.n163 AVSS.n162 0.0431396
R5178 AVSS.n162 AVSS.n161 0.0431396
R5179 AVSS.n73 AVSS.n72 0.0420736
R5180 AVSS.n428 AVSS.n427 0.041314
R5181 AVSS.n398 AVSS.n397 0.041314
R5182 AVSS.n273 AVSS.n272 0.041314
R5183 AVSS.n431 AVSS.n430 0.0411047
R5184 AVSS.n188 AVSS.n187 0.0411047
R5185 AVSS.n388 AVSS.n387 0.0411047
R5186 AVSS.n477 AVSS.n476 0.039811
R5187 AVSS.n269 AVSS.n268 0.039811
R5188 AVSS.n424 AVSS.n423 0.0385295
R5189 AVSS.n402 AVSS.n401 0.0385295
R5190 AVSS.n134 AVSS.n133 0.0365464
R5191 AVSS.n102 AVSS.n101 0.0364399
R5192 AVSS.n366 AVSS.n365 0.0354077
R5193 AVSS.n358 AVSS.n357 0.0354077
R5194 AVSS.n296 AVSS.n295 0.0354077
R5195 AVSS.n288 AVSS.n287 0.0354077
R5196 AVSS.n409 AVSS.n408 0.0353617
R5197 AVSS.n417 AVSS.n416 0.0353617
R5198 AVSS.n103 AVSS.n102 0.0346894
R5199 AVSS.n105 AVSS.n104 0.0346894
R5200 AVSS.n137 AVSS.n136 0.0346894
R5201 AVSS.n135 AVSS.n134 0.0346894
R5202 AVSS.n443 AVSS.n442 0.0342762
R5203 AVSS.n123 AVSS.n122 0.0342758
R5204 AVSS.n372 AVSS.n347 0.0337454
R5205 AVSS.n370 AVSS.n347 0.0337454
R5206 AVSS.n370 AVSS.n369 0.0337454
R5207 AVSS.n369 AVSS.n368 0.0337454
R5208 AVSS.n368 AVSS.n348 0.0337454
R5209 AVSS.n366 AVSS.n348 0.0337454
R5210 AVSS.n365 AVSS.n349 0.0337454
R5211 AVSS.n363 AVSS.n349 0.0337454
R5212 AVSS.n363 AVSS.n362 0.0337454
R5213 AVSS.n360 AVSS.n359 0.0337454
R5214 AVSS.n359 AVSS.n358 0.0337454
R5215 AVSS.n357 AVSS.n350 0.0337454
R5216 AVSS.n355 AVSS.n350 0.0337454
R5217 AVSS.n355 AVSS.n354 0.0337454
R5218 AVSS.n354 AVSS.n353 0.0337454
R5219 AVSS.n353 AVSS.n351 0.0337454
R5220 AVSS.n351 AVSS.n10 0.0337454
R5221 AVSS.n302 AVSS.n275 0.0337454
R5222 AVSS.n300 AVSS.n275 0.0337454
R5223 AVSS.n300 AVSS.n299 0.0337454
R5224 AVSS.n299 AVSS.n298 0.0337454
R5225 AVSS.n298 AVSS.n276 0.0337454
R5226 AVSS.n296 AVSS.n276 0.0337454
R5227 AVSS.n295 AVSS.n277 0.0337454
R5228 AVSS.n293 AVSS.n277 0.0337454
R5229 AVSS.n293 AVSS.n292 0.0337454
R5230 AVSS.n290 AVSS.n278 0.0337454
R5231 AVSS.n288 AVSS.n278 0.0337454
R5232 AVSS.n287 AVSS.n279 0.0337454
R5233 AVSS.n285 AVSS.n279 0.0337454
R5234 AVSS.n285 AVSS.n284 0.0337454
R5235 AVSS.n284 AVSS.n283 0.0337454
R5236 AVSS.n283 AVSS.n280 0.0337454
R5237 AVSS.n281 AVSS.n280 0.0337454
R5238 AVSS.n402 AVSS.n181 0.0337016
R5239 AVSS.n404 AVSS.n181 0.0337016
R5240 AVSS.n405 AVSS.n404 0.0337016
R5241 AVSS.n406 AVSS.n405 0.0337016
R5242 AVSS.n406 AVSS.n180 0.0337016
R5243 AVSS.n408 AVSS.n180 0.0337016
R5244 AVSS.n409 AVSS.n179 0.0337016
R5245 AVSS.n411 AVSS.n179 0.0337016
R5246 AVSS.n412 AVSS.n411 0.0337016
R5247 AVSS.n414 AVSS.n178 0.0337016
R5248 AVSS.n416 AVSS.n178 0.0337016
R5249 AVSS.n417 AVSS.n177 0.0337016
R5250 AVSS.n419 AVSS.n177 0.0337016
R5251 AVSS.n420 AVSS.n419 0.0337016
R5252 AVSS.n421 AVSS.n420 0.0337016
R5253 AVSS.n421 AVSS.n176 0.0337016
R5254 AVSS.n423 AVSS.n176 0.0337016
R5255 AVSS.n360 AVSS.n65 0.033033
R5256 AVSS.n291 AVSS.n290 0.033033
R5257 AVSS.n414 AVSS.n413 0.0329901
R5258 AVSS.n159 AVSS.n74 0.032073
R5259 AVSS.n124 AVSS.n123 0.0319607
R5260 AVSS.n125 AVSS.n124 0.0319607
R5261 AVSS.n125 AVSS.n110 0.0319607
R5262 AVSS.n127 AVSS.n110 0.0319607
R5263 AVSS.n130 AVSS.n129 0.0319607
R5264 AVSS.n131 AVSS.n130 0.0319607
R5265 AVSS.n131 AVSS.n109 0.0319607
R5266 AVSS.n133 AVSS.n109 0.0319607
R5267 AVSS.n92 AVSS.n74 0.0319607
R5268 AVSS.n93 AVSS.n92 0.0319607
R5269 AVSS.n93 AVSS.n91 0.0319607
R5270 AVSS.n95 AVSS.n91 0.0319607
R5271 AVSS.n98 AVSS.n97 0.0319607
R5272 AVSS.n99 AVSS.n98 0.0319607
R5273 AVSS.n99 AVSS.n90 0.0319607
R5274 AVSS.n101 AVSS.n90 0.0319607
R5275 AVSS.n202 AVSS.n60 0.0319161
R5276 AVSS.n484 AVSS.n483 0.0315563
R5277 AVSS.n262 AVSS.n261 0.0315563
R5278 AVSS.n476 AVSS.n475 0.0314767
R5279 AVSS.n425 AVSS.n424 0.0314767
R5280 AVSS.n427 AVSS.n426 0.0314767
R5281 AVSS.n429 AVSS.n428 0.0314767
R5282 AVSS.n432 AVSS.n431 0.0314767
R5283 AVSS.n430 AVSS.n0 0.0314767
R5284 AVSS.n401 AVSS.n400 0.0314767
R5285 AVSS.n399 AVSS.n398 0.0314767
R5286 AVSS.n397 AVSS.n396 0.0314767
R5287 AVSS.n187 AVSS.n182 0.0314767
R5288 AVSS.n189 AVSS.n188 0.0314767
R5289 AVSS.n270 AVSS.n269 0.0314767
R5290 AVSS.n272 AVSS.n271 0.0314767
R5291 AVSS.n274 AVSS.n273 0.0314767
R5292 AVSS.n389 AVSS.n388 0.0314767
R5293 AVSS.n387 AVSS.n386 0.0314767
R5294 AVSS.n385 AVSS.n384 0.0314767
R5295 AVSS.n486 AVSS.n485 0.0300775
R5296 AVSS.n485 AVSS.n484 0.0300775
R5297 AVSS.n483 AVSS.n4 0.0300775
R5298 AVSS.n481 AVSS.n4 0.0300775
R5299 AVSS.n481 AVSS.n480 0.0300775
R5300 AVSS.n480 AVSS.n479 0.0300775
R5301 AVSS.n479 AVSS.n5 0.0300775
R5302 AVSS.n477 AVSS.n5 0.0300775
R5303 AVSS.n268 AVSS.n183 0.0300775
R5304 AVSS.n266 AVSS.n183 0.0300775
R5305 AVSS.n266 AVSS.n265 0.0300775
R5306 AVSS.n265 AVSS.n264 0.0300775
R5307 AVSS.n264 AVSS.n184 0.0300775
R5308 AVSS.n262 AVSS.n184 0.0300775
R5309 AVSS.n261 AVSS.n185 0.0300775
R5310 AVSS.n259 AVSS.n185 0.0300775
R5311 AVSS.n259 AVSS.n258 0.0300775
R5312 AVSS.n161 AVSS.n160 0.0280818
R5313 AVSS.n472 AVSS.n9 0.0277138
R5314 AVSS.n471 AVSS.n10 0.0271502
R5315 AVSS.n166 AVSS.n165 0.0259315
R5316 AVSS.n115 AVSS.n114 0.0255699
R5317 AVSS.n486 AVSS.n3 0.0231186
R5318 AVSS.n474 AVSS.n473 0.0217442
R5319 AVSS.n384 AVSS.n383 0.0213083
R5320 AVSS.n204 AVSS.n203 0.0209545
R5321 AVSS.n445 AVSS.n444 0.0208496
R5322 AVSS.n373 AVSS.n372 0.0206172
R5323 AVSS.n383 AVSS.n302 0.0206172
R5324 AVSS.n281 AVSS.n58 0.0204409
R5325 AVSS.n138 AVSS.n137 0.0185
R5326 AVSS.n154 AVSS.n153 0.0181748
R5327 AVSS.n118 AVSS.n116 0.0173337
R5328 AVSS.n120 AVSS.n116 0.0173337
R5329 AVSS.n108 AVSS.n105 0.0172219
R5330 AVSS.n117 AVSS.n71 0.0169128
R5331 AVSS.n373 AVSS.n346 0.016599
R5332 AVSS.n122 AVSS.n121 0.0164441
R5333 AVSS.n112 AVSS.n111 0.0160769
R5334 AVSS.n205 AVSS.n204 0.0160245
R5335 AVSS.n203 AVSS.n202 0.0160245
R5336 AVSS.n444 AVSS.n443 0.0160245
R5337 AVSS.n446 AVSS.n445 0.0160245
R5338 AVSS.n346 AVSS.n58 0.0158871
R5339 AVSS.n257 AVSS.n256 0.0157873
R5340 AVSS.n129 AVSS.n128 0.0156685
R5341 AVSS.n97 AVSS.n96 0.0156685
R5342 AVSS.n472 AVSS.n471 0.0137679
R5343 AVSS.n128 AVSS.n127 0.0136461
R5344 AVSS.n96 AVSS.n95 0.0136461
R5345 AVSS.n155 AVSS.n154 0.0118287
R5346 AVSS.n157 AVSS.n156 0.011514
R5347 AVSS.n473 AVSS.n9 0.0113855
R5348 AVSS.n448 AVSS.n59 0.0113305
R5349 AVSS.n114 AVSS.n113 0.0105699
R5350 AVSS.n121 AVSS.n120 0.0105401
R5351 AVSS.n151 AVSS.n75 0.00999301
R5352 AVSS.n253 AVSS.n252 0.00799437
R5353 AVSS.n241 AVSS.n240 0.00799437
R5354 AVSS.n254 AVSS.n192 0.00752176
R5355 AVSS.n200 AVSS.n199 0.00752176
R5356 AVSS.n239 AVSS.n201 0.00752176
R5357 AVSS.n231 AVSS.n230 0.007488
R5358 AVSS.n219 AVSS.n218 0.007488
R5359 AVSS.n145 AVSS.n81 0.00721329
R5360 AVSS.n7 AVSS.n6 0.00704376
R5361 AVSS.n168 AVSS.n69 0.00704376
R5362 AVSS.n167 AVSS.n69 0.00704376
R5363 AVSS.n211 AVSS.n210 0.00701538
R5364 AVSS.n228 AVSS.n212 0.00701538
R5365 AVSS.n227 AVSS.n213 0.00701538
R5366 AVSS.n215 AVSS.n214 0.00701538
R5367 AVSS.n224 AVSS.n223 0.00701538
R5368 AVSS.n222 AVSS.n221 0.00701538
R5369 AVSS.n238 AVSS.n206 0.00684659
R5370 AVSS.n194 AVSS.n193 0.00667779
R5371 AVSS.n250 AVSS.n195 0.00667779
R5372 AVSS.n249 AVSS.n196 0.00667779
R5373 AVSS.n198 AVSS.n197 0.00667779
R5374 AVSS.n246 AVSS.n245 0.00667779
R5375 AVSS.n244 AVSS.n243 0.00667779
R5376 AVSS.n156 AVSS.n155 0.00653147
R5377 AVSS.n158 AVSS.n157 0.00632168
R5378 AVSS.n448 AVSS.n447 0.00619059
R5379 AVSS.n190 AVSS.n186 0.00617142
R5380 AVSS.n235 AVSS.n234 0.00617142
R5381 AVSS.n233 AVSS.n232 0.00617142
R5382 AVSS.n217 AVSS.n216 0.00617142
R5383 AVSS.n2 AVSS.n1 0.00617142
R5384 AVSS.n79 AVSS.n75 0.00611189
R5385 AVSS.n209 AVSS.n208 0.00596887
R5386 AVSS.n80 AVSS.n79 0.00490559
R5387 AVSS.n68 AVSS.n8 0.00489366
R5388 AVSS.n169 AVSS.n168 0.00489366
R5389 AVSS.n473 AVSS.n8 0.00442625
R5390 AVSS.n146 AVSS.n80 0.00432867
R5391 AVSS.n235 AVSS.n209 0.00428095
R5392 AVSS.n234 AVSS.n233 0.00428095
R5393 AVSS.n232 AVSS.n231 0.00428095
R5394 AVSS.n218 AVSS.n217 0.00428095
R5395 AVSS.n491 AVSS.n490 0.00428095
R5396 AVSS.n489 AVSS.n1 0.00428095
R5397 AVSS.n160 AVSS.n159 0.00385664
R5398 AVSS.n252 AVSS.n193 0.00377457
R5399 AVSS.n195 AVSS.n194 0.00377457
R5400 AVSS.n250 AVSS.n249 0.00377457
R5401 AVSS.n197 AVSS.n196 0.00377457
R5402 AVSS.n246 AVSS.n198 0.00377457
R5403 AVSS.n245 AVSS.n244 0.00377457
R5404 AVSS.n243 AVSS.n241 0.00377457
R5405 AVSS.n216 AVSS 0.00370705
R5406 AVSS.n207 AVSS.n206 0.00360578
R5407 AVSS.n230 AVSS.n210 0.00343698
R5408 AVSS.n212 AVSS.n211 0.00343698
R5409 AVSS.n228 AVSS.n227 0.00343698
R5410 AVSS.n214 AVSS.n213 0.00343698
R5411 AVSS.n224 AVSS.n215 0.00343698
R5412 AVSS.n223 AVSS.n222 0.00343698
R5413 AVSS.n221 AVSS.n219 0.00343698
R5414 AVSS.n473 AVSS.n6 0.0031175
R5415 AVSS.n442 AVSS.n60 0.00296504
R5416 AVSS.n256 AVSS.n186 0.00293061
R5417 AVSS.n192 AVSS.n191 0.00293061
R5418 AVSS.n254 AVSS.n253 0.00293061
R5419 AVSS.n240 AVSS.n199 0.00293061
R5420 AVSS.n201 AVSS.n200 0.00293061
R5421 AVSS.n239 AVSS.n238 0.00293061
R5422 AVSS.n346 AVSS.n59 0.00286014
R5423 AVSS.n159 AVSS.n158 0.00265035
R5424 AVSS.n111 AVSS.n81 0.00265035
R5425 AVSS.n490 AVSS.n489 0.00239047
R5426 AVSS.n152 AVSS.n151 0.00223077
R5427 AVSS.n138 AVSS.n108 0.00209763
R5428 AVSS.n191 AVSS.n190 0.00185034
R5429 AVSS.n113 AVSS.n112 0.00175874
R5430 AVSS.n313 AVSS.n310 0.00168421
R5431 AVSS.n377 AVSS.n308 0.00168421
R5432 AVSS.n380 AVSS.n305 0.00168421
R5433 AVSS.n468 AVSS.n467 0.00168421
R5434 AVSS.n464 AVSS.n463 0.00168421
R5435 AVSS.n459 AVSS.n458 0.00168421
R5436 AVSS.n455 AVSS.n454 0.00168421
R5437 AVSS.n31 AVSS.n30 0.00168421
R5438 AVSS.n27 AVSS.n26 0.00168421
R5439 AVSS.n22 AVSS.n21 0.00168421
R5440 AVSS.n140 AVSS.n88 0.00168421
R5441 AVSS.n143 AVSS.n84 0.00168421
R5442 AVSS.n163 AVSS.n73 0.00156599
R5443 AVSS.n167 AVSS.n166 0.00155167
R5444 AVSS.n121 AVSS.n115 0.00139161
R5445 AVSS.n146 AVSS.n145 0.00128671
R5446 AVSS.n362 AVSS.n65 0.0012124
R5447 AVSS.n292 AVSS.n291 0.0012124
R5448 AVSS.n413 AVSS.n412 0.00121146
R5449 AVSS.n258 AVSS.n257 0.0011338
R5450 AVSS.n491 AVSS 0.00107389
R5451 AVSS.n118 AVSS.n117 0.000920842
R5452 AVSS.n208 AVSS.n207 0.000702551
R5453 AVSS.n3 AVSS.n2 0.000702551
R5454 AVSS.n153 AVSS.n152 0.000604895
R5455 a_5396_n6451.t63 a_5396_n6451.t2 9.46371
R5456 a_5396_n6451.t16 a_5396_n6451.t52 8.7152
R5457 a_5396_n6451.t47 a_5396_n6451.t54 8.7152
R5458 a_5396_n6451.n7 a_5396_n6451.t156 9.1601
R5459 a_5396_n6451.n11 a_5396_n6451.t84 9.1601
R5460 a_5396_n6451.n25 a_5396_n6451.t88 9.17607
R5461 a_5396_n6451.n17 a_5396_n6451.t134 9.17607
R5462 a_5396_n6451.n110 a_5396_n6451.t140 8.10567
R5463 a_5396_n6451.n96 a_5396_n6451.t72 8.10567
R5464 a_5396_n6451.n96 a_5396_n6451.t164 8.10567
R5465 a_5396_n6451.n96 a_5396_n6451.t158 8.10567
R5466 a_5396_n6451.n96 a_5396_n6451.t211 8.10567
R5467 a_5396_n6451.n55 a_5396_n6451.t69 8.10567
R5468 a_5396_n6451.n55 a_5396_n6451.t236 8.10567
R5469 a_5396_n6451.n55 a_5396_n6451.t110 8.10567
R5470 a_5396_n6451.n55 a_5396_n6451.t100 8.10567
R5471 a_5396_n6451.n59 a_5396_n6451.t152 8.10567
R5472 a_5396_n6451.n59 a_5396_n6451.t206 8.10567
R5473 a_5396_n6451.n59 a_5396_n6451.t194 8.10567
R5474 a_5396_n6451.n59 a_5396_n6451.t71 8.10567
R5475 a_5396_n6451.n93 a_5396_n6451.t127 8.10567
R5476 a_5396_n6451.n93 a_5396_n6451.t118 8.10567
R5477 a_5396_n6451.n93 a_5396_n6451.t169 8.10567
R5478 a_5396_n6451.n91 a_5396_n6451.t212 8.10567
R5479 a_5396_n6451.n91 a_5396_n6451.t200 8.10567
R5480 a_5396_n6451.n91 a_5396_n6451.t79 8.10567
R5481 a_5396_n6451.n110 a_5396_n6451.t132 8.10567
R5482 a_5396_n6451.n110 a_5396_n6451.t209 8.10567
R5483 a_5396_n6451.n110 a_5396_n6451.t196 8.10567
R5484 a_5396_n6451.n116 a_5396_n6451.t198 8.10567
R5485 a_5396_n6451.n107 a_5396_n6451.t170 8.10567
R5486 a_5396_n6451.n107 a_5396_n6451.t231 8.10567
R5487 a_5396_n6451.n107 a_5396_n6451.t190 8.10567
R5488 a_5396_n6451.n107 a_5396_n6451.t133 8.10567
R5489 a_5396_n6451.n75 a_5396_n6451.t218 8.10567
R5490 a_5396_n6451.n75 a_5396_n6451.t175 8.10567
R5491 a_5396_n6451.n75 a_5396_n6451.t103 8.10567
R5492 a_5396_n6451.n75 a_5396_n6451.t240 8.10567
R5493 a_5396_n6451.n72 a_5396_n6451.t146 8.10567
R5494 a_5396_n6451.n72 a_5396_n6451.t90 8.10567
R5495 a_5396_n6451.n72 a_5396_n6451.t214 8.10567
R5496 a_5396_n6451.n72 a_5396_n6451.t149 8.10567
R5497 a_5396_n6451.n103 a_5396_n6451.t124 8.10567
R5498 a_5396_n6451.n103 a_5396_n6451.t87 8.10567
R5499 a_5396_n6451.n103 a_5396_n6451.t203 8.10567
R5500 a_5396_n6451.n78 a_5396_n6451.t97 8.10567
R5501 a_5396_n6451.n78 a_5396_n6451.t235 8.10567
R5502 a_5396_n6451.n78 a_5396_n6451.t177 8.10567
R5503 a_5396_n6451.n116 a_5396_n6451.t160 8.10567
R5504 a_5396_n6451.n116 a_5396_n6451.t119 8.10567
R5505 a_5396_n6451.n116 a_5396_n6451.t82 8.10567
R5506 a_5396_n6451.n112 a_5396_n6451.t187 8.10567
R5507 a_5396_n6451.n97 a_5396_n6451.t159 8.10567
R5508 a_5396_n6451.n97 a_5396_n6451.t222 8.10567
R5509 a_5396_n6451.n97 a_5396_n6451.t179 8.10567
R5510 a_5396_n6451.n97 a_5396_n6451.t122 8.10567
R5511 a_5396_n6451.n63 a_5396_n6451.t205 8.10567
R5512 a_5396_n6451.n63 a_5396_n6451.t165 8.10567
R5513 a_5396_n6451.n63 a_5396_n6451.t94 8.10567
R5514 a_5396_n6451.n63 a_5396_n6451.t232 8.10567
R5515 a_5396_n6451.n68 a_5396_n6451.t135 8.10567
R5516 a_5396_n6451.n68 a_5396_n6451.t80 8.10567
R5517 a_5396_n6451.n68 a_5396_n6451.t197 8.10567
R5518 a_5396_n6451.n68 a_5396_n6451.t142 8.10567
R5519 a_5396_n6451.n89 a_5396_n6451.t99 8.10567
R5520 a_5396_n6451.n89 a_5396_n6451.t239 8.10567
R5521 a_5396_n6451.n89 a_5396_n6451.t181 8.10567
R5522 a_5396_n6451.n66 a_5396_n6451.t78 8.10567
R5523 a_5396_n6451.n66 a_5396_n6451.t215 8.10567
R5524 a_5396_n6451.n66 a_5396_n6451.t154 8.10567
R5525 a_5396_n6451.n112 a_5396_n6451.t148 8.10567
R5526 a_5396_n6451.n112 a_5396_n6451.t108 8.10567
R5527 a_5396_n6451.n112 a_5396_n6451.t70 8.10567
R5528 a_5396_n6451.n115 a_5396_n6451.t126 8.10567
R5529 a_5396_n6451.n106 a_5396_n6451.t96 8.10567
R5530 a_5396_n6451.n106 a_5396_n6451.t157 8.10567
R5531 a_5396_n6451.n106 a_5396_n6451.t117 8.10567
R5532 a_5396_n6451.n106 a_5396_n6451.t234 8.10567
R5533 a_5396_n6451.n85 a_5396_n6451.t143 8.10567
R5534 a_5396_n6451.n85 a_5396_n6451.t106 8.10567
R5535 a_5396_n6451.n85 a_5396_n6451.t207 8.10567
R5536 a_5396_n6451.n85 a_5396_n6451.t166 8.10567
R5537 a_5396_n6451.n86 a_5396_n6451.t75 8.10567
R5538 a_5396_n6451.n86 a_5396_n6451.t189 8.10567
R5539 a_5396_n6451.n86 a_5396_n6451.t137 8.10567
R5540 a_5396_n6451.n86 a_5396_n6451.t81 8.10567
R5541 a_5396_n6451.n101 a_5396_n6451.t230 8.10567
R5542 a_5396_n6451.n101 a_5396_n6451.t186 8.10567
R5543 a_5396_n6451.n101 a_5396_n6451.t130 8.10567
R5544 a_5396_n6451.n99 a_5396_n6451.t201 8.10567
R5545 a_5396_n6451.n99 a_5396_n6451.t163 8.10567
R5546 a_5396_n6451.n99 a_5396_n6451.t107 8.10567
R5547 a_5396_n6451.n115 a_5396_n6451.t91 8.10567
R5548 a_5396_n6451.n115 a_5396_n6451.t225 8.10567
R5549 a_5396_n6451.n115 a_5396_n6451.t183 8.10567
R5550 a_5396_n6451.n13 a_5396_n6451.t85 8.10567
R5551 a_5396_n6451.n13 a_5396_n6451.t77 8.10567
R5552 a_5396_n6451.n13 a_5396_n6451.t125 8.10567
R5553 a_5396_n6451.n13 a_5396_n6451.t115 8.10567
R5554 a_5396_n6451.n165 a_5396_n6451.t112 8.10567
R5555 a_5396_n6451.n166 a_5396_n6451.t102 8.10567
R5556 a_5396_n6451.n12 a_5396_n6451.t153 8.10567
R5557 a_5396_n6451.n26 a_5396_n6451.t180 8.10567
R5558 a_5396_n6451.n26 a_5396_n6451.t171 8.10567
R5559 a_5396_n6451.n26 a_5396_n6451.t227 8.10567
R5560 a_5396_n6451.n2 a_5396_n6451.t155 8.10567
R5561 a_5396_n6451.n2 a_5396_n6451.t147 8.10567
R5562 a_5396_n6451.n2 a_5396_n6451.t226 8.10567
R5563 a_5396_n6451.n39 a_5396_n6451.t193 8.10567
R5564 a_5396_n6451.n146 a_5396_n6451.t185 8.10567
R5565 a_5396_n6451.n145 a_5396_n6451.t237 8.10567
R5566 a_5396_n6451.n40 a_5396_n6451.t168 8.10567
R5567 a_5396_n6451.n40 a_5396_n6451.t223 8.10567
R5568 a_5396_n6451.n41 a_5396_n6451.t213 8.10567
R5569 a_5396_n6451.n41 a_5396_n6451.t86 8.10567
R5570 a_5396_n6451.n36 a_5396_n6451.t199 8.10567
R5571 a_5396_n6451.n36 a_5396_n6451.t161 8.10567
R5572 a_5396_n6451.n36 a_5396_n6451.t89 8.10567
R5573 a_5396_n6451.n36 a_5396_n6451.t228 8.10567
R5574 a_5396_n6451.n149 a_5396_n6451.t139 8.10567
R5575 a_5396_n6451.n150 a_5396_n6451.t98 8.10567
R5576 a_5396_n6451.n35 a_5396_n6451.t220 8.10567
R5577 a_5396_n6451.n8 a_5396_n6451.t217 8.10567
R5578 a_5396_n6451.n8 a_5396_n6451.t174 8.10567
R5579 a_5396_n6451.n8 a_5396_n6451.t116 8.10567
R5580 a_5396_n6451.n29 a_5396_n6451.t184 8.10567
R5581 a_5396_n6451.n29 a_5396_n6451.t145 8.10567
R5582 a_5396_n6451.n29 a_5396_n6451.t105 8.10567
R5583 a_5396_n6451.n50 a_5396_n6451.t114 8.10567
R5584 a_5396_n6451.n148 a_5396_n6451.t76 8.10567
R5585 a_5396_n6451.n147 a_5396_n6451.t192 8.10567
R5586 a_5396_n6451.n46 a_5396_n6451.t131 8.10567
R5587 a_5396_n6451.n46 a_5396_n6451.t73 8.10567
R5588 a_5396_n6451.n51 a_5396_n6451.t195 8.10567
R5589 a_5396_n6451.n51 a_5396_n6451.t136 8.10567
R5590 a_5396_n6451.n23 a_5396_n6451.t176 8.10567
R5591 a_5396_n6451.n23 a_5396_n6451.t138 8.10567
R5592 a_5396_n6451.n23 a_5396_n6451.t67 8.10567
R5593 a_5396_n6451.n23 a_5396_n6451.t202 8.10567
R5594 a_5396_n6451.n15 a_5396_n6451.t129 8.10567
R5595 a_5396_n6451.n156 a_5396_n6451.t93 8.10567
R5596 a_5396_n6451.n155 a_5396_n6451.t210 8.10567
R5597 a_5396_n6451.n16 a_5396_n6451.t191 8.10567
R5598 a_5396_n6451.n16 a_5396_n6451.t151 8.10567
R5599 a_5396_n6451.n16 a_5396_n6451.t95 8.10567
R5600 a_5396_n6451.n4 a_5396_n6451.t162 8.10567
R5601 a_5396_n6451.n4 a_5396_n6451.t123 8.10567
R5602 a_5396_n6451.n4 a_5396_n6451.t83 8.10567
R5603 a_5396_n6451.n37 a_5396_n6451.t104 8.10567
R5604 a_5396_n6451.n154 a_5396_n6451.t241 8.10567
R5605 a_5396_n6451.n153 a_5396_n6451.t182 8.10567
R5606 a_5396_n6451.n20 a_5396_n6451.t109 8.10567
R5607 a_5396_n6451.n20 a_5396_n6451.t229 8.10567
R5608 a_5396_n6451.n38 a_5396_n6451.t172 8.10567
R5609 a_5396_n6451.n38 a_5396_n6451.t113 8.10567
R5610 a_5396_n6451.n34 a_5396_n6451.t128 8.10567
R5611 a_5396_n6451.n34 a_5396_n6451.t92 8.10567
R5612 a_5396_n6451.n34 a_5396_n6451.t188 8.10567
R5613 a_5396_n6451.n34 a_5396_n6451.t150 8.10567
R5614 a_5396_n6451.n9 a_5396_n6451.t68 8.10567
R5615 a_5396_n6451.n162 a_5396_n6451.t204 8.10567
R5616 a_5396_n6451.n161 a_5396_n6451.t144 8.10567
R5617 a_5396_n6451.n10 a_5396_n6451.t141 8.10567
R5618 a_5396_n6451.n10 a_5396_n6451.t101 8.10567
R5619 a_5396_n6451.n10 a_5396_n6451.t224 8.10567
R5620 a_5396_n6451.n31 a_5396_n6451.t111 8.10567
R5621 a_5396_n6451.n31 a_5396_n6451.t74 8.10567
R5622 a_5396_n6451.n31 a_5396_n6451.t208 8.10567
R5623 a_5396_n6451.n48 a_5396_n6451.t219 8.10567
R5624 a_5396_n6451.n160 a_5396_n6451.t178 8.10567
R5625 a_5396_n6451.n159 a_5396_n6451.t120 8.10567
R5626 a_5396_n6451.n43 a_5396_n6451.t233 8.10567
R5627 a_5396_n6451.n43 a_5396_n6451.t173 8.10567
R5628 a_5396_n6451.n45 a_5396_n6451.t121 8.10567
R5629 a_5396_n6451.n45 a_5396_n6451.t238 8.10567
R5630 a_5396_n6451.t25 a_5396_n6451.t16 7.22198
R5631 a_5396_n6451.t21 a_5396_n6451.t47 7.22198
R5632 a_5396_n6451.t1 a_5396_n6451.t4 7.12006
R5633 a_5396_n6451.n187 a_5396_n6451.t11 6.77653
R5634 a_5396_n6451.n177 a_5396_n6451.t41 6.77653
R5635 a_5396_n6451.n190 a_5396_n6451.t56 6.7761
R5636 a_5396_n6451.t5 a_5396_n6451.n216 6.7761
R5637 a_5396_n6451.n138 a_5396_n6451.t66 6.86989
R5638 a_5396_n6451.n127 a_5396_n6451.t62 6.77231
R5639 a_5396_n6451.n137 a_5396_n6451.t15 6.77231
R5640 a_5396_n6451.n194 a_5396_n6451.t3 6.14835
R5641 a_5396_n6451.n192 a_5396_n6451.t65 6.14517
R5642 a_5396_n6451.t10 a_5396_n6451.t9 5.70489
R5643 a_5396_n6451.t30 a_5396_n6451.t31 5.70489
R5644 a_5396_n6451.n191 a_5396_n6451.t64 5.61877
R5645 a_5396_n6451.n139 a_5396_n6451.t8 5.50607
R5646 a_5396_n6451.n178 a_5396_n6451.t59 5.50607
R5647 a_5396_n6451.n205 a_5396_n6451.t42 5.50607
R5648 a_5396_n6451.n188 a_5396_n6451.t23 5.50607
R5649 a_5396_n6451.n177 a_5396_n6451.t18 5.50475
R5650 a_5396_n6451.n180 a_5396_n6451.t12 5.50475
R5651 a_5396_n6451.n183 a_5396_n6451.t20 5.50475
R5652 a_5396_n6451.n187 a_5396_n6451.t39 5.50475
R5653 a_5396_n6451.n190 a_5396_n6451.t24 5.50475
R5654 a_5396_n6451.n206 a_5396_n6451.t51 5.50475
R5655 a_5396_n6451.n209 a_5396_n6451.t7 5.50475
R5656 a_5396_n6451.n216 a_5396_n6451.t28 5.50475
R5657 a_5396_n6451.n181 a_5396_n6451.t37 5.50475
R5658 a_5396_n6451.n182 a_5396_n6451.t55 5.50475
R5659 a_5396_n6451.n179 a_5396_n6451.t6 5.50475
R5660 a_5396_n6451.n204 a_5396_n6451.t34 5.50475
R5661 a_5396_n6451.n207 a_5396_n6451.t45 5.50475
R5662 a_5396_n6451.n208 a_5396_n6451.t29 5.50475
R5663 a_5396_n6451.n189 a_5396_n6451.t61 5.50475
R5664 a_5396_n6451.n88 a_5396_n6451.n40 0.595624
R5665 a_5396_n6451.n21 a_5396_n6451.n20 0.595624
R5666 a_5396_n6451.n47 a_5396_n6451.n46 0.607617
R5667 a_5396_n6451.n32 a_5396_n6451.n43 0.607617
R5668 a_5396_n6451.n118 a_5396_n6451.t14 5.5012
R5669 a_5396_n6451.n119 a_5396_n6451.t46 5.5012
R5670 a_5396_n6451.n120 a_5396_n6451.t49 5.5012
R5671 a_5396_n6451.n121 a_5396_n6451.t26 5.5012
R5672 a_5396_n6451.n122 a_5396_n6451.t38 5.5012
R5673 a_5396_n6451.n123 a_5396_n6451.t33 5.5012
R5674 a_5396_n6451.n124 a_5396_n6451.t44 5.5012
R5675 a_5396_n6451.t58 a_5396_n6451.n125 5.5012
R5676 a_5396_n6451.t60 a_5396_n6451.n126 5.5012
R5677 a_5396_n6451.t53 a_5396_n6451.n127 5.5012
R5678 a_5396_n6451.n128 a_5396_n6451.t22 5.5012
R5679 a_5396_n6451.t50 a_5396_n6451.n129 5.5012
R5680 a_5396_n6451.t27 a_5396_n6451.n130 5.5012
R5681 a_5396_n6451.t13 a_5396_n6451.n131 5.5012
R5682 a_5396_n6451.t43 a_5396_n6451.n132 5.5012
R5683 a_5396_n6451.t40 a_5396_n6451.n133 5.5012
R5684 a_5396_n6451.t48 a_5396_n6451.n134 5.5012
R5685 a_5396_n6451.t36 a_5396_n6451.n135 5.5012
R5686 a_5396_n6451.t57 a_5396_n6451.n136 5.5012
R5687 a_5396_n6451.t35 a_5396_n6451.n137 5.5012
R5688 a_5396_n6451.t0 a_5396_n6451.n138 5.66099
R5689 a_5396_n6451.n108 a_5396_n6451.n107 0.020246
R5690 a_5396_n6451.n106 a_5396_n6451.n105 0.020246
R5691 a_5396_n6451.n75 a_5396_n6451.n74 0.150803
R5692 a_5396_n6451.n73 a_5396_n6451.n72 0.150806
R5693 a_5396_n6451.n116 a_5396_n6451.n77 0.0676355
R5694 a_5396_n6451.n85 a_5396_n6451.n83 0.150783
R5695 a_5396_n6451.n86 a_5396_n6451.n82 0.150803
R5696 a_5396_n6451.n115 a_5396_n6451.n114 0.0676355
R5697 a_5396_n6451.n60 a_5396_n6451.n59 0.153625
R5698 a_5396_n6451.n56 a_5396_n6451.n55 0.153625
R5699 a_5396_n6451.n96 a_5396_n6451.n95 0.020088
R5700 a_5396_n6451.n72 a_5396_n6451.n80 0.246907
R5701 a_5396_n6451.n76 a_5396_n6451.n75 0.246907
R5702 a_5396_n6451.n68 a_5396_n6451.n61 0.153625
R5703 a_5396_n6451.n63 a_5396_n6451.n62 0.153625
R5704 a_5396_n6451.n98 a_5396_n6451.n97 0.020088
R5705 a_5396_n6451.n112 a_5396_n6451.n65 0.0201939
R5706 a_5396_n6451.n69 a_5396_n6451.n68 0.246907
R5707 a_5396_n6451.n64 a_5396_n6451.n63 0.246907
R5708 a_5396_n6451.n87 a_5396_n6451.n86 0.246907
R5709 a_5396_n6451.n85 a_5396_n6451.n84 0.246877
R5710 a_5396_n6451.n110 a_5396_n6451.n109 0.0201939
R5711 a_5396_n6451.n59 a_5396_n6451.n58 0.246907
R5712 a_5396_n6451.n55 a_5396_n6451.n54 0.246907
R5713 a_5396_n6451.n29 a_5396_n6451.n28 0.260442
R5714 a_5396_n6451.n52 a_5396_n6451.n51 0.591264
R5715 a_5396_n6451.n36 a_5396_n6451.n5 0.310971
R5716 a_5396_n6451.n8 a_5396_n6451.n7 0.258567
R5717 a_5396_n6451.n4 a_5396_n6451.n3 0.208479
R5718 a_5396_n6451.n38 a_5396_n6451.n19 0.591642
R5719 a_5396_n6451.n23 a_5396_n6451.n22 0.623337
R5720 a_5396_n6451.n17 a_5396_n6451.n16 0.259585
R5721 a_5396_n6451.n31 a_5396_n6451.n30 0.260442
R5722 a_5396_n6451.n49 a_5396_n6451.n45 0.591264
R5723 a_5396_n6451.n34 a_5396_n6451.n33 0.310971
R5724 a_5396_n6451.n11 a_5396_n6451.n10 0.258567
R5725 a_5396_n6451.n2 a_5396_n6451.n1 0.208479
R5726 a_5396_n6451.n42 a_5396_n6451.n41 0.591642
R5727 a_5396_n6451.n14 a_5396_n6451.n13 0.623337
R5728 a_5396_n6451.n26 a_5396_n6451.n25 0.259585
R5729 a_5396_n6451.n200 a_5396_n6451.n196 3.48654
R5730 a_5396_n6451.n197 a_5396_n6451.n196 3.42822
R5731 a_5396_n6451.n176 a_5396_n6451.n175 3.37173
R5732 a_5396_n6451.n139 a_5396_n6451.t17 3.32015
R5733 a_5396_n6451.n215 a_5396_n6451.t30 3.23904
R5734 a_5396_n6451.n201 a_5396_n6451.t10 3.23904
R5735 a_5396_n6451.n193 a_5396_n6451.t1 3.23004
R5736 a_5396_n6451.n208 a_5396_n6451.n207 2.60203
R5737 a_5396_n6451.n182 a_5396_n6451.n181 2.60203
R5738 a_5396_n6451.n189 a_5396_n6451.n188 2.52436
R5739 a_5396_n6451.n205 a_5396_n6451.n204 2.52436
R5740 a_5396_n6451.n179 a_5396_n6451.n178 2.52436
R5741 a_5396_n6451.n173 a_5396_n6451.n168 2.40699
R5742 a_5396_n6451.n151 a_5396_n6451.n27 2.30989
R5743 a_5396_n6451.n157 a_5396_n6451.n6 2.30989
R5744 a_5396_n6451.n193 a_5396_n6451.n192 2.2807
R5745 a_5396_n6451.n94 a_5396_n6451.n93 0.427602
R5746 a_5396_n6451.n92 a_5396_n6451.n91 0.427602
R5747 a_5396_n6451.n90 a_5396_n6451.n89 0.427602
R5748 a_5396_n6451.n67 a_5396_n6451.n66 0.427602
R5749 a_5396_n6451.n104 a_5396_n6451.n103 0.420727
R5750 a_5396_n6451.n79 a_5396_n6451.n78 0.420727
R5751 a_5396_n6451.n102 a_5396_n6451.n101 0.420727
R5752 a_5396_n6451.n100 a_5396_n6451.n99 0.420727
R5753 a_5396_n6451.n111 a_5396_n6451.n69 2.96488
R5754 a_5396_n6451.n98 a_5396_n6451.n117 2.94096
R5755 a_5396_n6451.n58 a_5396_n6451.n57 2.96488
R5756 a_5396_n6451.n53 a_5396_n6451.n95 2.94096
R5757 a_5396_n6451.n171 a_5396_n6451.n71 2.07182
R5758 a_5396_n6451.n170 a_5396_n6451.n70 2.07182
R5759 a_5396_n6451.n73 a_5396_n6451.n71 2.75704
R5760 a_5396_n6451.n70 a_5396_n6451.n108 2.90773
R5761 a_5396_n6451.n113 a_5396_n6451.n82 2.75706
R5762 a_5396_n6451.n105 a_5396_n6451.n81 2.90773
R5763 a_5396_n6451.n175 a_5396_n6451.n174 1.80314
R5764 a_5396_n6451.n140 a_5396_n6451.n141 1.70908
R5765 a_5396_n6451.n168 a_5396_n6451.n167 1.68395
R5766 a_5396_n6451.n164 a_5396_n6451.n141 1.68395
R5767 a_5396_n6451.n172 a_5396_n6451.n113 1.5005
R5768 a_5396_n6451.n171 a_5396_n6451.n111 1.5005
R5769 a_5396_n6451.n57 a_5396_n6451.n173 1.5005
R5770 a_5396_n6451.n174 a_5396_n6451.n53 1.5005
R5771 a_5396_n6451.n81 a_5396_n6451.n169 1.5005
R5772 a_5396_n6451.n117 a_5396_n6451.n170 1.5005
R5773 a_5396_n6451.n158 a_5396_n6451.n144 1.5005
R5774 a_5396_n6451.n152 a_5396_n6451.n151 1.5005
R5775 a_5396_n6451.n167 a_5396_n6451.n0 1.5005
R5776 a_5396_n6451.n24 a_5396_n6451.n164 1.5005
R5777 a_5396_n6451.n163 a_5396_n6451.n44 1.5005
R5778 a_5396_n6451.n157 a_5396_n6451.n18 1.5005
R5779 a_5396_n6451.n198 a_5396_n6451.n197 1.5005
R5780 a_5396_n6451.t47 a_5396_n6451.n186 1.5005
R5781 a_5396_n6451.n211 a_5396_n6451.n210 1.5005
R5782 a_5396_n6451.n214 a_5396_n6451.n213 1.5005
R5783 a_5396_n6451.t16 a_5396_n6451.n143 1.5005
R5784 a_5396_n6451.n195 a_5396_n6451.n194 1.5005
R5785 a_5396_n6451.n200 a_5396_n6451.n199 1.5005
R5786 a_5396_n6451.n203 a_5396_n6451.n202 1.5005
R5787 a_5396_n6451.n212 a_5396_n6451.n142 1.5005
R5788 a_5396_n6451.t17 a_5396_n6451.n140 1.5005
R5789 a_5396_n6451.n185 a_5396_n6451.n184 1.5005
R5790 a_5396_n6451.n172 a_5396_n6451.n171 1.47516
R5791 a_5396_n6451.n170 a_5396_n6451.n169 1.47516
R5792 a_5396_n6451.n196 a_5396_n6451.n195 1.41182
R5793 a_5396_n6451.n28 a_5396_n6451.t242 9.17619
R5794 a_5396_n6451.n30 a_5396_n6451.t167 9.17619
R5795 a_5396_n6451.t30 a_5396_n6451.t25 1.27228
R5796 a_5396_n6451.n209 a_5396_n6451.n208 1.27228
R5797 a_5396_n6451.n207 a_5396_n6451.n206 1.27228
R5798 a_5396_n6451.t10 a_5396_n6451.t21 1.27228
R5799 a_5396_n6451.n183 a_5396_n6451.n182 1.27228
R5800 a_5396_n6451.n181 a_5396_n6451.n180 1.27228
R5801 a_5396_n6451.n188 a_5396_n6451.n187 1.26756
R5802 a_5396_n6451.n206 a_5396_n6451.n205 1.26756
R5803 a_5396_n6451.n178 a_5396_n6451.n177 1.26756
R5804 a_5396_n6451.n180 a_5396_n6451.n139 1.26756
R5805 a_5396_n6451.n149 a_5396_n6451.n8 1.24866
R5806 a_5396_n6451.n51 a_5396_n6451.n50 1.24866
R5807 a_5396_n6451.n10 a_5396_n6451.n9 1.24866
R5808 a_5396_n6451.n45 a_5396_n6451.n48 1.24866
R5809 a_5396_n6451.n147 a_5396_n6451.n29 1.24629
R5810 a_5396_n6451.n159 a_5396_n6451.n31 1.24629
R5811 a_5396_n6451.n151 a_5396_n6451.n144 1.23709
R5812 a_5396_n6451.n163 a_5396_n6451.n157 1.23709
R5813 a_5396_n6451.n13 a_5396_n6451.n12 1.22261
R5814 a_5396_n6451.n145 a_5396_n6451.n2 1.22261
R5815 a_5396_n6451.n155 a_5396_n6451.n23 1.22261
R5816 a_5396_n6451.n153 a_5396_n6451.n4 1.22261
R5817 a_5396_n6451.n165 a_5396_n6451.n26 1.21313
R5818 a_5396_n6451.n41 a_5396_n6451.n39 1.21313
R5819 a_5396_n6451.n16 a_5396_n6451.n15 1.21313
R5820 a_5396_n6451.n38 a_5396_n6451.n37 1.21313
R5821 a_5396_n6451.n185 a_5396_n6451.n176 1.10472
R5822 a_5396_n6451.n167 a_5396_n6451.n144 0.809892
R5823 a_5396_n6451.n164 a_5396_n6451.n163 0.809892
R5824 a_5396_n6451.n210 a_5396_n6451.n189 0.796291
R5825 a_5396_n6451.n204 a_5396_n6451.n203 0.796291
R5826 a_5396_n6451.n184 a_5396_n6451.n179 0.796291
R5827 a_5396_n6451.n143 a_5396_n6451.n214 0.780703
R5828 a_5396_n6451.n197 a_5396_n6451.n186 0.780703
R5829 a_5396_n6451.n215 a_5396_n6451.n142 0.780703
R5830 a_5396_n6451.n201 a_5396_n6451.n200 0.780703
R5831 a_5396_n6451.n194 a_5396_n6451.t63 0.769291
R5832 a_5396_n6451.n192 a_5396_n6451.n191 0.767125
R5833 a_5396_n6451.n27 a_5396_n6451.n52 1.14908
R5834 a_5396_n6451.n7 a_5396_n6451.n6 1.39299
R5835 a_5396_n6451.n49 a_5396_n6451.n158 1.14908
R5836 a_5396_n6451.n44 a_5396_n6451.n11 1.39299
R5837 a_5396_n6451.n152 a_5396_n6451.n19 1.11421
R5838 a_5396_n6451.n18 a_5396_n6451.n17 1.35707
R5839 a_5396_n6451.n0 a_5396_n6451.n42 1.11421
R5840 a_5396_n6451.n25 a_5396_n6451.n24 1.35707
R5841 a_5396_n6451.n12 a_5396_n6451.n166 0.673132
R5842 a_5396_n6451.n166 a_5396_n6451.n165 0.673132
R5843 a_5396_n6451.n146 a_5396_n6451.n145 0.673132
R5844 a_5396_n6451.n39 a_5396_n6451.n146 0.673132
R5845 a_5396_n6451.n35 a_5396_n6451.n150 0.673132
R5846 a_5396_n6451.n150 a_5396_n6451.n149 0.673132
R5847 a_5396_n6451.n148 a_5396_n6451.n147 0.673132
R5848 a_5396_n6451.n50 a_5396_n6451.n148 0.673132
R5849 a_5396_n6451.n156 a_5396_n6451.n155 0.673132
R5850 a_5396_n6451.n15 a_5396_n6451.n156 0.673132
R5851 a_5396_n6451.n154 a_5396_n6451.n153 0.673132
R5852 a_5396_n6451.n37 a_5396_n6451.n154 0.673132
R5853 a_5396_n6451.n162 a_5396_n6451.n161 0.673132
R5854 a_5396_n6451.n9 a_5396_n6451.n162 0.673132
R5855 a_5396_n6451.n160 a_5396_n6451.n159 0.673132
R5856 a_5396_n6451.n48 a_5396_n6451.n160 0.673132
R5857 a_5396_n6451.n143 a_5396_n6451.n185 0.638405
R5858 a_5396_n6451.n211 a_5396_n6451.n186 0.638405
R5859 a_5396_n6451.n195 a_5396_n6451.n193 0.638405
R5860 a_5396_n6451.n140 a_5396_n6451.n215 0.638405
R5861 a_5396_n6451.n202 a_5396_n6451.n201 0.638405
R5862 a_5396_n6451.n214 a_5396_n6451.n211 0.628372
R5863 a_5396_n6451.n202 a_5396_n6451.n142 0.628372
R5864 a_5396_n6451.n175 a_5396_n6451.n141 0.604355
R5865 a_5396_n6451.n176 a_5396_n6451.n168 0.603852
R5866 a_5396_n6451.n173 a_5396_n6451.n172 0.571818
R5867 a_5396_n6451.n174 a_5396_n6451.n169 0.571818
R5868 a_5396_n6451.n210 a_5396_n6451.n209 0.476484
R5869 a_5396_n6451.n203 a_5396_n6451.n190 0.476484
R5870 a_5396_n6451.n184 a_5396_n6451.n183 0.476484
R5871 a_5396_n6451.n216 a_5396_n6451.t17 0.476484
R5872 a_5396_n6451.n47 a_5396_n6451.n52 1.14166
R5873 a_5396_n6451.n6 a_5396_n6451.n5 2.75347
R5874 a_5396_n6451.n49 a_5396_n6451.n32 1.14166
R5875 a_5396_n6451.n44 a_5396_n6451.n33 2.75347
R5876 a_5396_n6451.n213 a_5396_n6451.n124 0.478684
R5877 a_5396_n6451.n212 a_5396_n6451.n118 0.478684
R5878 a_5396_n6451.n134 a_5396_n6451.n198 0.478684
R5879 a_5396_n6451.n199 a_5396_n6451.n128 0.478684
R5880 a_5396_n6451.n92 a_5396_n6451.n109 2.03311
R5881 a_5396_n6451.n60 a_5396_n6451.n92 2.04491
R5882 a_5396_n6451.n56 a_5396_n6451.n60 4.37762
R5883 a_5396_n6451.n94 a_5396_n6451.n56 1.87961
R5884 a_5396_n6451.n95 a_5396_n6451.n94 2.19836
R5885 a_5396_n6451.n79 a_5396_n6451.n77 2.03667
R5886 a_5396_n6451.n80 a_5396_n6451.n79 2.21715
R5887 a_5396_n6451.n76 a_5396_n6451.n80 4.49317
R5888 a_5396_n6451.n104 a_5396_n6451.n76 1.82113
R5889 a_5396_n6451.n108 a_5396_n6451.n104 2.19319
R5890 a_5396_n6451.n71 a_5396_n6451.n77 1.65342
R5891 a_5396_n6451.n74 a_5396_n6451.n73 4.34574
R5892 a_5396_n6451.n74 a_5396_n6451.n70 1.50586
R5893 a_5396_n6451.n67 a_5396_n6451.n65 2.03311
R5894 a_5396_n6451.n61 a_5396_n6451.n67 2.04491
R5895 a_5396_n6451.n62 a_5396_n6451.n61 4.37762
R5896 a_5396_n6451.n90 a_5396_n6451.n62 1.87961
R5897 a_5396_n6451.n90 a_5396_n6451.n98 2.19836
R5898 a_5396_n6451.n65 a_5396_n6451.n111 1.65903
R5899 a_5396_n6451.n69 a_5396_n6451.n64 4.49309
R5900 a_5396_n6451.n64 a_5396_n6451.n117 1.44546
R5901 a_5396_n6451.n100 a_5396_n6451.n114 2.03667
R5902 a_5396_n6451.n87 a_5396_n6451.n100 2.2172
R5903 a_5396_n6451.n87 a_5396_n6451.n84 4.49278
R5904 a_5396_n6451.n102 a_5396_n6451.n84 1.82125
R5905 a_5396_n6451.n102 a_5396_n6451.n105 2.19319
R5906 a_5396_n6451.n114 a_5396_n6451.n113 1.65342
R5907 a_5396_n6451.n83 a_5396_n6451.n82 4.34534
R5908 a_5396_n6451.n83 a_5396_n6451.n81 1.50598
R5909 a_5396_n6451.n57 a_5396_n6451.n109 1.65903
R5910 a_5396_n6451.n58 a_5396_n6451.n54 4.49309
R5911 a_5396_n6451.n54 a_5396_n6451.n53 1.44546
R5912 a_5396_n6451.n28 a_5396_n6451.n27 2.8103
R5913 a_5396_n6451.n47 a_5396_n6451.n5 4.38327
R5914 a_5396_n6451.n152 a_5396_n6451.n3 2.83621
R5915 a_5396_n6451.n21 a_5396_n6451.n19 1.15119
R5916 a_5396_n6451.n22 a_5396_n6451.n21 4.37089
R5917 a_5396_n6451.n22 a_5396_n6451.n18 2.6764
R5918 a_5396_n6451.n158 a_5396_n6451.n30 2.8103
R5919 a_5396_n6451.n33 a_5396_n6451.n32 4.38327
R5920 a_5396_n6451.n1 a_5396_n6451.n0 2.83621
R5921 a_5396_n6451.n42 a_5396_n6451.n88 1.15119
R5922 a_5396_n6451.n88 a_5396_n6451.n14 4.37089
R5923 a_5396_n6451.n14 a_5396_n6451.n24 2.6764
R5924 a_5396_n6451.n126 a_5396_n6451.n127 1.27228
R5925 a_5396_n6451.n125 a_5396_n6451.n126 2.51878
R5926 a_5396_n6451.n213 a_5396_n6451.n125 0.794091
R5927 a_5396_n6451.n123 a_5396_n6451.n124 1.27228
R5928 a_5396_n6451.n122 a_5396_n6451.n123 2.60203
R5929 a_5396_n6451.n121 a_5396_n6451.n122 1.27228
R5930 a_5396_n6451.n120 a_5396_n6451.n121 1.27228
R5931 a_5396_n6451.n119 a_5396_n6451.n120 2.51878
R5932 a_5396_n6451.n212 a_5396_n6451.n119 0.794091
R5933 a_5396_n6451.t19 a_5396_n6451.n118 6.77266
R5934 a_5396_n6451.n136 a_5396_n6451.n137 1.27228
R5935 a_5396_n6451.n135 a_5396_n6451.n136 2.51878
R5936 a_5396_n6451.n198 a_5396_n6451.n135 0.794091
R5937 a_5396_n6451.n133 a_5396_n6451.n134 1.27228
R5938 a_5396_n6451.n132 a_5396_n6451.n133 2.60203
R5939 a_5396_n6451.n131 a_5396_n6451.n132 1.27228
R5940 a_5396_n6451.n130 a_5396_n6451.n131 1.27228
R5941 a_5396_n6451.n129 a_5396_n6451.n130 2.51878
R5942 a_5396_n6451.n199 a_5396_n6451.n129 0.794091
R5943 a_5396_n6451.t32 a_5396_n6451.n128 6.77266
R5944 a_5396_n6451.n191 a_5396_n6451.n138 3.17898
R5945 a_5396_n6451.n41 a_5396_n6451.n40 2.16997
R5946 a_5396_n6451.n20 a_5396_n6451.n38 2.16997
R5947 a_5396_n6451.n36 a_5396_n6451.n35 2.13563
R5948 a_5396_n6451.n161 a_5396_n6451.n34 2.13563
R5949 a_5396_n6451.n51 a_5396_n6451.n46 2.13445
R5950 a_5396_n6451.n43 a_5396_n6451.n45 2.13445
R5951 a_5396_n6451.t221 a_5396_n6451.n3 9.16748
R5952 a_5396_n6451.t216 a_5396_n6451.n1 9.16748
R5953 a_5396_8177.n68 a_5396_8177.n67 7.22198
R5954 a_5396_8177.n179 a_5396_8177.n178 7.22198
R5955 a_5396_8177.n42 a_5396_8177.t0 6.77653
R5956 a_5396_8177.n38 a_5396_8177.t38 6.77653
R5957 a_5396_8177.n46 a_5396_8177.t41 6.7761
R5958 a_5396_8177.n192 a_5396_8177.t80 6.7761
R5959 a_5396_8177.n8 a_5396_8177.t11 6.77231
R5960 a_5396_8177.n18 a_5396_8177.t15 6.77231
R5961 a_5396_8177.n150 a_5396_8177.n149 6.50088
R5962 a_5396_8177.n115 a_5396_8177.n111 6.50088
R5963 a_5396_8177.n49 a_5396_8177.t21 5.50607
R5964 a_5396_8177.n43 a_5396_8177.t28 5.50607
R5965 a_5396_8177.n189 a_5396_8177.t56 5.50607
R5966 a_5396_8177.n39 a_5396_8177.t66 5.50607
R5967 a_5396_8177.n48 a_5396_8177.t61 5.50475
R5968 a_5396_8177.n52 a_5396_8177.t6 5.50475
R5969 a_5396_8177.n53 a_5396_8177.t54 5.50475
R5970 a_5396_8177.n44 a_5396_8177.t52 5.50475
R5971 a_5396_8177.n190 a_5396_8177.t9 5.50475
R5972 a_5396_8177.n186 a_5396_8177.t45 5.50475
R5973 a_5396_8177.n185 a_5396_8177.t4 5.50475
R5974 a_5396_8177.n40 a_5396_8177.t2 5.50475
R5975 a_5396_8177.n82 a_5396_8177.n80 4.92758
R5976 a_5396_8177.n121 a_5396_8177.n119 4.92758
R5977 a_5396_8177.n25 a_5396_8177.n88 4.92217
R5978 a_5396_8177.n32 a_5396_8177.n101 4.92217
R5979 a_5396_8177.n19 a_5396_8177.n95 3.65107
R5980 a_5396_8177.n20 a_5396_8177.n94 3.65107
R5981 a_5396_8177.n21 a_5396_8177.n93 3.65107
R5982 a_5396_8177.n22 a_5396_8177.n92 3.65107
R5983 a_5396_8177.n91 a_5396_8177.n23 3.65107
R5984 a_5396_8177.n90 a_5396_8177.n24 3.65107
R5985 a_5396_8177.n89 a_5396_8177.n25 3.65107
R5986 a_5396_8177.n26 a_5396_8177.n108 3.65107
R5987 a_5396_8177.n27 a_5396_8177.n107 3.65107
R5988 a_5396_8177.n28 a_5396_8177.n106 3.65107
R5989 a_5396_8177.n29 a_5396_8177.n105 3.65107
R5990 a_5396_8177.n104 a_5396_8177.n30 3.65107
R5991 a_5396_8177.n103 a_5396_8177.n31 3.65107
R5992 a_5396_8177.n102 a_5396_8177.n32 3.65107
R5993 a_5396_8177.n33 a_5396_8177.n197 4.0312
R5994 a_5396_8177.n0 a_5396_8177.n34 4.0312
R5995 a_5396_8177.n1 a_5396_8177.t73 5.5012
R5996 a_5396_8177.n2 a_5396_8177.t32 5.5012
R5997 a_5396_8177.n3 a_5396_8177.t20 5.5012
R5998 a_5396_8177.n4 a_5396_8177.t67 5.5012
R5999 a_5396_8177.n5 a_5396_8177.n71 4.0312
R6000 a_5396_8177.t64 a_5396_8177.n6 5.5012
R6001 a_5396_8177.t39 a_5396_8177.n7 5.5012
R6002 a_5396_8177.n70 a_5396_8177.n8 4.0312
R6003 a_5396_8177.n9 a_5396_8177.n78 4.0312
R6004 a_5396_8177.n10 a_5396_8177.t7 5.5012
R6005 a_5396_8177.n11 a_5396_8177.t79 5.5012
R6006 a_5396_8177.n12 a_5396_8177.n77 4.0312
R6007 a_5396_8177.n13 a_5396_8177.t62 5.5012
R6008 a_5396_8177.n14 a_5396_8177.t37 5.5012
R6009 a_5396_8177.n15 a_5396_8177.n76 4.0312
R6010 a_5396_8177.t78 a_5396_8177.n16 5.5012
R6011 a_5396_8177.t42 a_5396_8177.n17 5.5012
R6012 a_5396_8177.n75 a_5396_8177.n18 4.0312
R6013 a_5396_8177.n66 a_5396_8177.t17 4.24002
R6014 a_5396_8177.n57 a_5396_8177.t29 4.24002
R6015 a_5396_8177.n177 a_5396_8177.t43 4.24002
R6016 a_5396_8177.n168 a_5396_8177.t3 4.24002
R6017 a_5396_8177.n116 a_5396_8177.t134 4.06712
R6018 a_5396_8177.n99 a_5396_8177.t143 4.06712
R6019 a_5396_8177.n144 a_5396_8177.t124 4.06712
R6020 a_5396_8177.n142 a_5396_8177.t166 4.06712
R6021 a_5396_8177.n46 a_5396_8177.n45 4.03475
R6022 a_5396_8177.n51 a_5396_8177.n50 4.03475
R6023 a_5396_8177.n55 a_5396_8177.n54 4.03475
R6024 a_5396_8177.n42 a_5396_8177.n41 4.03475
R6025 a_5396_8177.n192 a_5396_8177.n191 4.03475
R6026 a_5396_8177.n188 a_5396_8177.n187 4.03475
R6027 a_5396_8177.n184 a_5396_8177.n183 4.03475
R6028 a_5396_8177.n38 a_5396_8177.n37 4.03475
R6029 a_5396_8177.n163 a_5396_8177.n74 3.97307
R6030 a_5396_8177.n145 a_5396_8177.n79 3.96014
R6031 a_5396_8177.n118 a_5396_8177.n117 3.96014
R6032 a_5396_8177.n116 a_5396_8177.t133 3.86107
R6033 a_5396_8177.n99 a_5396_8177.t142 3.86107
R6034 a_5396_8177.n144 a_5396_8177.t125 3.86107
R6035 a_5396_8177.n142 a_5396_8177.t168 3.86107
R6036 a_5396_8177.n84 a_5396_8177.n82 3.79678
R6037 a_5396_8177.n159 a_5396_8177.n157 3.79678
R6038 a_5396_8177.n123 a_5396_8177.n121 3.79678
R6039 a_5396_8177.n132 a_5396_8177.n130 3.79678
R6040 a_5396_8177.n66 a_5396_8177.t12 3.68818
R6041 a_5396_8177.n57 a_5396_8177.t24 3.68818
R6042 a_5396_8177.n177 a_5396_8177.t48 3.68818
R6043 a_5396_8177.n168 a_5396_8177.t60 3.68818
R6044 a_5396_8177.n161 a_5396_8177.n160 3.65581
R6045 a_5396_8177.n159 a_5396_8177.n158 3.65581
R6046 a_5396_8177.n157 a_5396_8177.n156 3.65581
R6047 a_5396_8177.n155 a_5396_8177.n154 3.65581
R6048 a_5396_8177.n86 a_5396_8177.n85 3.65581
R6049 a_5396_8177.n84 a_5396_8177.n83 3.65581
R6050 a_5396_8177.n82 a_5396_8177.n81 3.65581
R6051 a_5396_8177.n134 a_5396_8177.n133 3.65581
R6052 a_5396_8177.n132 a_5396_8177.n131 3.65581
R6053 a_5396_8177.n130 a_5396_8177.n129 3.65581
R6054 a_5396_8177.n128 a_5396_8177.n127 3.65581
R6055 a_5396_8177.n125 a_5396_8177.n124 3.65581
R6056 a_5396_8177.n123 a_5396_8177.n122 3.65581
R6057 a_5396_8177.n121 a_5396_8177.n120 3.65581
R6058 a_5396_8177.n155 a_5396_8177.n153 3.64443
R6059 a_5396_8177.n128 a_5396_8177.n126 3.64443
R6060 a_5396_8177.n137 a_5396_8177.n22 3.64223
R6061 a_5396_8177.n109 a_5396_8177.n29 3.64223
R6062 a_5396_8177.n65 a_5396_8177.n35 3.23904
R6063 a_5396_8177.n176 a_5396_8177.n36 3.23904
R6064 a_5396_8177.n64 a_5396_8177.n63 2.77002
R6065 a_5396_8177.n60 a_5396_8177.n59 2.77002
R6066 a_5396_8177.n175 a_5396_8177.n174 2.77002
R6067 a_5396_8177.n171 a_5396_8177.n170 2.77002
R6068 a_5396_8177.n61 a_5396_8177.n57 2.73714
R6069 a_5396_8177.n172 a_5396_8177.n168 2.73714
R6070 a_5396_8177.n143 a_5396_8177.n141 2.73714
R6071 a_5396_8177.n100 a_5396_8177.n98 2.73714
R6072 a_5396_8177.n53 a_5396_8177.n52 2.60203
R6073 a_5396_8177.n186 a_5396_8177.n185 2.60203
R6074 a_5396_8177.n114 a_5396_8177.n112 2.59712
R6075 a_5396_8177.n98 a_5396_8177.n96 2.59712
R6076 a_5396_8177.n148 a_5396_8177.n146 2.59712
R6077 a_5396_8177.n141 a_5396_8177.n139 2.59712
R6078 a_5396_8177.n44 a_5396_8177.n43 2.52436
R6079 a_5396_8177.n49 a_5396_8177.n48 2.52436
R6080 a_5396_8177.n40 a_5396_8177.n39 2.52436
R6081 a_5396_8177.n190 a_5396_8177.n189 2.52436
R6082 a_5396_8177.n150 a_5396_8177.n143 2.46014
R6083 a_5396_8177.n111 a_5396_8177.n100 2.46014
R6084 a_5396_8177.n114 a_5396_8177.n113 2.39107
R6085 a_5396_8177.n98 a_5396_8177.n97 2.39107
R6086 a_5396_8177.n148 a_5396_8177.n147 2.39107
R6087 a_5396_8177.n141 a_5396_8177.n140 2.39107
R6088 a_5396_8177.n64 a_5396_8177.n62 2.21818
R6089 a_5396_8177.n60 a_5396_8177.n58 2.21818
R6090 a_5396_8177.n175 a_5396_8177.n173 2.21818
R6091 a_5396_8177.n171 a_5396_8177.n169 2.21818
R6092 a_5396_8177.n69 a_5396_8177.n56 2.13841
R6093 a_5396_8177.n47 a_5396_8177.n35 2.13841
R6094 a_5396_8177.n110 a_5396_8177.n109 2.0852
R6095 a_5396_8177.n163 a_5396_8177.n162 2.02864
R6096 a_5396_8177.n167 a_5396_8177.n74 1.76168
R6097 a_5396_8177.n68 a_5396_8177.n61 1.73904
R6098 a_5396_8177.n179 a_5396_8177.n172 1.73904
R6099 a_5396_8177.n162 a_5396_8177.n161 1.73609
R6100 a_5396_8177.n135 a_5396_8177.n134 1.73609
R6101 a_5396_8177.n167 a_5396_8177.n166 1.5005
R6102 a_5396_8177.n180 a_5396_8177.n179 1.5005
R6103 a_5396_8177.n182 a_5396_8177.n181 1.5005
R6104 a_5396_8177.n69 a_5396_8177.n68 1.5005
R6105 a_5396_8177.n151 a_5396_8177.n150 1.5005
R6106 a_5396_8177.n126 a_5396_8177.n87 1.5005
R6107 a_5396_8177.n138 a_5396_8177.n137 1.5005
R6108 a_5396_8177.n153 a_5396_8177.n152 1.5005
R6109 a_5396_8177.n111 a_5396_8177.n110 1.5005
R6110 a_5396_8177.n165 a_5396_8177.n164 1.5005
R6111 a_5396_8177.n194 a_5396_8177.n193 1.5005
R6112 a_5396_8177.n196 a_5396_8177.n195 1.5005
R6113 a_5396_8177.n73 a_5396_8177.n72 1.5005
R6114 a_5396_8177.n34 a_5396_8177.t44 1.4705
R6115 a_5396_8177.n34 a_5396_8177.t25 1.4705
R6116 a_5396_8177.n71 a_5396_8177.t35 1.4705
R6117 a_5396_8177.n71 a_5396_8177.t5 1.4705
R6118 a_5396_8177.n70 a_5396_8177.t81 1.4705
R6119 a_5396_8177.n70 a_5396_8177.t58 1.4705
R6120 a_5396_8177.n45 a_5396_8177.t33 1.4705
R6121 a_5396_8177.n45 a_5396_8177.t14 1.4705
R6122 a_5396_8177.n50 a_5396_8177.t76 1.4705
R6123 a_5396_8177.n50 a_5396_8177.t40 1.4705
R6124 a_5396_8177.n54 a_5396_8177.t22 1.4705
R6125 a_5396_8177.n54 a_5396_8177.t85 1.4705
R6126 a_5396_8177.n41 a_5396_8177.t68 1.4705
R6127 a_5396_8177.n41 a_5396_8177.t47 1.4705
R6128 a_5396_8177.n62 a_5396_8177.t72 1.4705
R6129 a_5396_8177.n62 a_5396_8177.t50 1.4705
R6130 a_5396_8177.n63 a_5396_8177.t74 1.4705
R6131 a_5396_8177.n63 a_5396_8177.t55 1.4705
R6132 a_5396_8177.n58 a_5396_8177.t83 1.4705
R6133 a_5396_8177.n58 a_5396_8177.t63 1.4705
R6134 a_5396_8177.n59 a_5396_8177.t1 1.4705
R6135 a_5396_8177.n59 a_5396_8177.t69 1.4705
R6136 a_5396_8177.n191 a_5396_8177.t71 1.4705
R6137 a_5396_8177.n191 a_5396_8177.t49 1.4705
R6138 a_5396_8177.n187 a_5396_8177.t26 1.4705
R6139 a_5396_8177.n187 a_5396_8177.t75 1.4705
R6140 a_5396_8177.n183 a_5396_8177.t59 1.4705
R6141 a_5396_8177.n183 a_5396_8177.t34 1.4705
R6142 a_5396_8177.n37 a_5396_8177.t18 1.4705
R6143 a_5396_8177.n37 a_5396_8177.t84 1.4705
R6144 a_5396_8177.n173 a_5396_8177.t19 1.4705
R6145 a_5396_8177.n173 a_5396_8177.t86 1.4705
R6146 a_5396_8177.n174 a_5396_8177.t70 1.4705
R6147 a_5396_8177.n174 a_5396_8177.t65 1.4705
R6148 a_5396_8177.n169 a_5396_8177.t31 1.4705
R6149 a_5396_8177.n169 a_5396_8177.t13 1.4705
R6150 a_5396_8177.n170 a_5396_8177.t27 1.4705
R6151 a_5396_8177.n170 a_5396_8177.t23 1.4705
R6152 a_5396_8177.n78 a_5396_8177.t36 1.4705
R6153 a_5396_8177.n78 a_5396_8177.t30 1.4705
R6154 a_5396_8177.n77 a_5396_8177.t57 1.4705
R6155 a_5396_8177.n77 a_5396_8177.t82 1.4705
R6156 a_5396_8177.n76 a_5396_8177.t16 1.4705
R6157 a_5396_8177.n76 a_5396_8177.t10 1.4705
R6158 a_5396_8177.n75 a_5396_8177.t8 1.4705
R6159 a_5396_8177.n75 a_5396_8177.t46 1.4705
R6160 a_5396_8177.n112 a_5396_8177.t95 1.4705
R6161 a_5396_8177.n112 a_5396_8177.t154 1.4705
R6162 a_5396_8177.n113 a_5396_8177.t93 1.4705
R6163 a_5396_8177.n113 a_5396_8177.t153 1.4705
R6164 a_5396_8177.n96 a_5396_8177.t106 1.4705
R6165 a_5396_8177.n96 a_5396_8177.t162 1.4705
R6166 a_5396_8177.n97 a_5396_8177.t105 1.4705
R6167 a_5396_8177.n97 a_5396_8177.t161 1.4705
R6168 a_5396_8177.n160 a_5396_8177.t103 1.4705
R6169 a_5396_8177.n160 a_5396_8177.t149 1.4705
R6170 a_5396_8177.n158 a_5396_8177.t169 1.4705
R6171 a_5396_8177.n158 a_5396_8177.t109 1.4705
R6172 a_5396_8177.n156 a_5396_8177.t156 1.4705
R6173 a_5396_8177.n156 a_5396_8177.t152 1.4705
R6174 a_5396_8177.n154 a_5396_8177.t136 1.4705
R6175 a_5396_8177.n154 a_5396_8177.t132 1.4705
R6176 a_5396_8177.n85 a_5396_8177.t172 1.4705
R6177 a_5396_8177.n85 a_5396_8177.t110 1.4705
R6178 a_5396_8177.n83 a_5396_8177.t150 1.4705
R6179 a_5396_8177.n83 a_5396_8177.t90 1.4705
R6180 a_5396_8177.n81 a_5396_8177.t121 1.4705
R6181 a_5396_8177.n81 a_5396_8177.t118 1.4705
R6182 a_5396_8177.n80 a_5396_8177.t88 1.4705
R6183 a_5396_8177.n80 a_5396_8177.t170 1.4705
R6184 a_5396_8177.n95 a_5396_8177.t158 1.4705
R6185 a_5396_8177.n95 a_5396_8177.t171 1.4705
R6186 a_5396_8177.n94 a_5396_8177.t160 1.4705
R6187 a_5396_8177.n94 a_5396_8177.t108 1.4705
R6188 a_5396_8177.n93 a_5396_8177.t115 1.4705
R6189 a_5396_8177.n93 a_5396_8177.t164 1.4705
R6190 a_5396_8177.n92 a_5396_8177.t137 1.4705
R6191 a_5396_8177.n92 a_5396_8177.t100 1.4705
R6192 a_5396_8177.n91 a_5396_8177.t94 1.4705
R6193 a_5396_8177.n91 a_5396_8177.t127 1.4705
R6194 a_5396_8177.n90 a_5396_8177.t116 1.4705
R6195 a_5396_8177.n90 a_5396_8177.t144 1.4705
R6196 a_5396_8177.n89 a_5396_8177.t148 1.4705
R6197 a_5396_8177.n89 a_5396_8177.t119 1.4705
R6198 a_5396_8177.n88 a_5396_8177.t175 1.4705
R6199 a_5396_8177.n88 a_5396_8177.t113 1.4705
R6200 a_5396_8177.n133 a_5396_8177.t165 1.4705
R6201 a_5396_8177.n133 a_5396_8177.t111 1.4705
R6202 a_5396_8177.n131 a_5396_8177.t130 1.4705
R6203 a_5396_8177.n131 a_5396_8177.t98 1.4705
R6204 a_5396_8177.n129 a_5396_8177.t107 1.4705
R6205 a_5396_8177.n129 a_5396_8177.t89 1.4705
R6206 a_5396_8177.n127 a_5396_8177.t159 1.4705
R6207 a_5396_8177.n127 a_5396_8177.t141 1.4705
R6208 a_5396_8177.n124 a_5396_8177.t151 1.4705
R6209 a_5396_8177.n124 a_5396_8177.t123 1.4705
R6210 a_5396_8177.n122 a_5396_8177.t120 1.4705
R6211 a_5396_8177.n122 a_5396_8177.t92 1.4705
R6212 a_5396_8177.n120 a_5396_8177.t117 1.4705
R6213 a_5396_8177.n120 a_5396_8177.t97 1.4705
R6214 a_5396_8177.n119 a_5396_8177.t155 1.4705
R6215 a_5396_8177.n119 a_5396_8177.t138 1.4705
R6216 a_5396_8177.n108 a_5396_8177.t96 1.4705
R6217 a_5396_8177.n108 a_5396_8177.t126 1.4705
R6218 a_5396_8177.n107 a_5396_8177.t140 1.4705
R6219 a_5396_8177.n107 a_5396_8177.t114 1.4705
R6220 a_5396_8177.n106 a_5396_8177.t122 1.4705
R6221 a_5396_8177.n106 a_5396_8177.t101 1.4705
R6222 a_5396_8177.n105 a_5396_8177.t91 1.4705
R6223 a_5396_8177.n105 a_5396_8177.t157 1.4705
R6224 a_5396_8177.n104 a_5396_8177.t163 1.4705
R6225 a_5396_8177.n104 a_5396_8177.t139 1.4705
R6226 a_5396_8177.n103 a_5396_8177.t135 1.4705
R6227 a_5396_8177.n103 a_5396_8177.t104 1.4705
R6228 a_5396_8177.n102 a_5396_8177.t131 1.4705
R6229 a_5396_8177.n102 a_5396_8177.t112 1.4705
R6230 a_5396_8177.n101 a_5396_8177.t167 1.4705
R6231 a_5396_8177.n101 a_5396_8177.t147 1.4705
R6232 a_5396_8177.n146 a_5396_8177.t99 1.4705
R6233 a_5396_8177.n146 a_5396_8177.t128 1.4705
R6234 a_5396_8177.n147 a_5396_8177.t102 1.4705
R6235 a_5396_8177.n147 a_5396_8177.t129 1.4705
R6236 a_5396_8177.n139 a_5396_8177.t145 1.4705
R6237 a_5396_8177.n139 a_5396_8177.t173 1.4705
R6238 a_5396_8177.n140 a_5396_8177.t146 1.4705
R6239 a_5396_8177.n140 a_5396_8177.t174 1.4705
R6240 a_5396_8177.t87 a_5396_8177.n197 1.4705
R6241 a_5396_8177.n197 a_5396_8177.t51 1.4705
R6242 a_5396_8177.n65 a_5396_8177.n64 1.46537
R6243 a_5396_8177.n67 a_5396_8177.n66 1.46537
R6244 a_5396_8177.n61 a_5396_8177.n60 1.46537
R6245 a_5396_8177.n176 a_5396_8177.n175 1.46537
R6246 a_5396_8177.n178 a_5396_8177.n177 1.46537
R6247 a_5396_8177.n172 a_5396_8177.n171 1.46537
R6248 a_5396_8177.n117 a_5396_8177.n116 1.46537
R6249 a_5396_8177.n115 a_5396_8177.n114 1.46537
R6250 a_5396_8177.n100 a_5396_8177.n99 1.46537
R6251 a_5396_8177.n145 a_5396_8177.n144 1.46537
R6252 a_5396_8177.n149 a_5396_8177.n148 1.46537
R6253 a_5396_8177.n143 a_5396_8177.n142 1.46537
R6254 a_5396_8177.n152 a_5396_8177.n74 1.42428
R6255 a_5396_8177.n55 a_5396_8177.n53 1.27228
R6256 a_5396_8177.n52 a_5396_8177.n51 1.27228
R6257 a_5396_8177.n67 a_5396_8177.n65 1.27228
R6258 a_5396_8177.n185 a_5396_8177.n184 1.27228
R6259 a_5396_8177.n188 a_5396_8177.n186 1.27228
R6260 a_5396_8177.n178 a_5396_8177.n176 1.27228
R6261 a_5396_8177.n86 a_5396_8177.n84 1.27228
R6262 a_5396_8177.n157 a_5396_8177.n155 1.27228
R6263 a_5396_8177.n161 a_5396_8177.n159 1.27228
R6264 a_5396_8177.n125 a_5396_8177.n123 1.27228
R6265 a_5396_8177.n130 a_5396_8177.n128 1.27228
R6266 a_5396_8177.n134 a_5396_8177.n132 1.27228
R6267 a_5396_8177.n149 a_5396_8177.n145 1.27228
R6268 a_5396_8177.n117 a_5396_8177.n115 1.27228
R6269 a_5396_8177.n43 a_5396_8177.n42 1.26756
R6270 a_5396_8177.n51 a_5396_8177.n49 1.26756
R6271 a_5396_8177.n39 a_5396_8177.n38 1.26756
R6272 a_5396_8177.n189 a_5396_8177.n188 1.26756
R6273 a_5396_8177.n164 a_5396_8177.n163 1.15732
R6274 a_5396_8177.n138 a_5396_8177.n87 0.822966
R6275 a_5396_8177.n136 a_5396_8177.n135 0.822966
R6276 a_5396_8177.n56 a_5396_8177.n44 0.796291
R6277 a_5396_8177.n48 a_5396_8177.n47 0.796291
R6278 a_5396_8177.n182 a_5396_8177.n40 0.796291
R6279 a_5396_8177.n193 a_5396_8177.n190 0.796291
R6280 a_5396_8177.n73 a_5396_8177.n69 0.780703
R6281 a_5396_8177.n180 a_5396_8177.n167 0.780703
R6282 a_5396_8177.n195 a_5396_8177.n35 0.780703
R6283 a_5396_8177.n164 a_5396_8177.n36 0.780703
R6284 a_5396_8177.n152 a_5396_8177.n151 0.639318
R6285 a_5396_8177.n110 a_5396_8177.n87 0.639318
R6286 a_5396_8177.n162 a_5396_8177.n79 0.639318
R6287 a_5396_8177.n135 a_5396_8177.n118 0.639318
R6288 a_5396_8177.n181 a_5396_8177.n180 0.638405
R6289 a_5396_8177.n194 a_5396_8177.n36 0.638405
R6290 a_5396_8177.n181 a_5396_8177.n73 0.628372
R6291 a_5396_8177.n195 a_5396_8177.n194 0.628372
R6292 a_5396_8177.n151 a_5396_8177.n138 0.585196
R6293 a_5396_8177.n136 a_5396_8177.n79 0.585196
R6294 a_5396_8177.n56 a_5396_8177.n55 0.476484
R6295 a_5396_8177.n47 a_5396_8177.n46 0.476484
R6296 a_5396_8177.n184 a_5396_8177.n182 0.476484
R6297 a_5396_8177.n193 a_5396_8177.n192 0.476484
R6298 a_5396_8177.n166 a_5396_8177.n15 0.478684
R6299 a_5396_8177.n165 a_5396_8177.n9 0.478684
R6300 a_5396_8177.n72 a_5396_8177.n5 0.478684
R6301 a_5396_8177.n196 a_5396_8177.n0 0.478684
R6302 a_5396_8177.n153 a_5396_8177.n86 0.236091
R6303 a_5396_8177.n126 a_5396_8177.n125 0.236091
R6304 a_5396_8177.n17 a_5396_8177.n18 1.27228
R6305 a_5396_8177.n16 a_5396_8177.n17 2.51878
R6306 a_5396_8177.n166 a_5396_8177.n16 0.794091
R6307 a_5396_8177.n14 a_5396_8177.n15 1.27228
R6308 a_5396_8177.n13 a_5396_8177.n14 2.60203
R6309 a_5396_8177.n12 a_5396_8177.n13 1.27228
R6310 a_5396_8177.n11 a_5396_8177.n12 1.27228
R6311 a_5396_8177.n10 a_5396_8177.n11 2.51878
R6312 a_5396_8177.n165 a_5396_8177.n10 0.794091
R6313 a_5396_8177.t77 a_5396_8177.n9 6.77266
R6314 a_5396_8177.n24 a_5396_8177.n25 3.79678
R6315 a_5396_8177.n23 a_5396_8177.n24 1.27228
R6316 a_5396_8177.n137 a_5396_8177.n23 0.238291
R6317 a_5396_8177.n21 a_5396_8177.n22 1.27228
R6318 a_5396_8177.n20 a_5396_8177.n21 3.79678
R6319 a_5396_8177.n19 a_5396_8177.n20 1.27228
R6320 a_5396_8177.n136 a_5396_8177.n19 1.73829
R6321 a_5396_8177.n31 a_5396_8177.n32 3.79678
R6322 a_5396_8177.n30 a_5396_8177.n31 1.27228
R6323 a_5396_8177.n109 a_5396_8177.n30 0.238291
R6324 a_5396_8177.n28 a_5396_8177.n29 1.27228
R6325 a_5396_8177.n27 a_5396_8177.n28 3.79678
R6326 a_5396_8177.n26 a_5396_8177.n27 1.27228
R6327 a_5396_8177.n26 a_5396_8177.n118 2.32299
R6328 a_5396_8177.n7 a_5396_8177.n8 1.27228
R6329 a_5396_8177.n6 a_5396_8177.n7 2.51878
R6330 a_5396_8177.n72 a_5396_8177.n6 0.794091
R6331 a_5396_8177.n4 a_5396_8177.n5 1.27228
R6332 a_5396_8177.n3 a_5396_8177.n4 2.60203
R6333 a_5396_8177.n33 a_5396_8177.n3 1.27263
R6334 a_5396_8177.n33 a_5396_8177.n2 1.27192
R6335 a_5396_8177.n1 a_5396_8177.n2 2.51878
R6336 a_5396_8177.n196 a_5396_8177.n1 0.794091
R6337 a_5396_8177.t53 a_5396_8177.n0 6.77266
R6338 IREF.n1383 IREF.n1292 16.7377
R6339 IREF.n1293 IREF.t22 10.214
R6340 IREF.n1303 IREF.t50 10.214
R6341 IREF.n1314 IREF.t179 10.214
R6342 IREF.n1325 IREF.t106 10.214
R6343 IREF.n1336 IREF.t181 10.214
R6344 IREF.n1299 IREF.t8 10.2117
R6345 IREF.n1309 IREF.t141 10.2117
R6346 IREF.n1320 IREF.t55 10.2117
R6347 IREF.n1331 IREF.t203 10.2117
R6348 IREF.n1342 IREF.t57 10.2117
R6349 IREF.n1296 IREF.t211 9.58832
R6350 IREF.n1306 IREF.t118 9.58832
R6351 IREF.n1317 IREF.t2 9.58832
R6352 IREF.n1364 IREF.t234 9.58832
R6353 IREF.n1328 IREF.t16 9.58832
R6354 IREF.n1339 IREF.t250 9.58832
R6355 IREF.n1298 IREF.t249 9.58085
R6356 IREF.n1308 IREF.t168 9.58085
R6357 IREF.n1319 IREF.t34 9.58085
R6358 IREF.n1366 IREF.t68 9.58085
R6359 IREF.n1330 IREF.t6 9.58085
R6360 IREF.n1341 IREF.t89 9.58085
R6361 IREF.n1297 IREF.t241 9.58045
R6362 IREF.n1295 IREF.t28 9.58045
R6363 IREF.n1294 IREF.t40 9.58045
R6364 IREF.n1307 IREF.t159 9.58045
R6365 IREF.n1305 IREF.t233 9.58045
R6366 IREF.n1304 IREF.t201 9.58045
R6367 IREF.n1318 IREF.t38 9.58045
R6368 IREF.n1316 IREF.t145 9.58045
R6369 IREF.n1315 IREF.t107 9.58045
R6370 IREF.n1365 IREF.t54 9.58045
R6371 IREF.n1329 IREF.t12 9.58045
R6372 IREF.n1327 IREF.t81 9.58045
R6373 IREF.n1326 IREF.t253 9.58045
R6374 IREF.n1340 IREF.t80 9.58045
R6375 IREF.n1338 IREF.t149 9.58045
R6376 IREF.n1337 IREF.t108 9.58045
R6377 IREF.n1293 IREF.t42 9.58005
R6378 IREF.n1303 IREF.t187 9.58005
R6379 IREF.n1314 IREF.t97 9.58005
R6380 IREF.n1325 IREF.t243 9.58005
R6381 IREF.n1336 IREF.t100 9.58005
R6382 IREF.n1299 IREF.t32 9.57886
R6383 IREF.n1300 IREF.t20 9.57886
R6384 IREF.n1301 IREF.t10 9.57886
R6385 IREF.n1309 IREF.t228 9.57886
R6386 IREF.n1310 IREF.t76 9.57886
R6387 IREF.n1311 IREF.t130 9.57886
R6388 IREF.n1320 IREF.t133 9.57886
R6389 IREF.n1321 IREF.t202 9.57886
R6390 IREF.n1322 IREF.t261 9.57886
R6391 IREF.n1331 IREF.t66 9.57886
R6392 IREF.n1332 IREF.t121 9.57886
R6393 IREF.n1333 IREF.t192 9.57886
R6394 IREF.n1342 IREF.t134 9.57886
R6395 IREF.n1343 IREF.t205 9.57886
R6396 IREF.n1344 IREF.t44 9.57886
R6397 IREF.n1370 IREF.t0 8.38951
R6398 IREF.n1351 IREF.t18 8.38752
R6399 IREF.n823 IREF.t176 8.38704
R6400 IREF.n805 IREF.t160 8.38704
R6401 IREF.n937 IREF.t46 8.37857
R6402 IREF.n1060 IREF.t173 8.37857
R6403 IREF.n870 IREF.t207 8.31301
R6404 IREF.n1021 IREF.t111 8.31301
R6405 IREF.n1170 IREF.t254 8.29322
R6406 IREF.n959 IREF.t237 8.29322
R6407 IREF.n80 IREF.t245 8.10567
R6408 IREF.n1213 IREF.t235 8.10567
R6409 IREF.n1207 IREF.t93 8.10567
R6410 IREF.n1202 IREF.t185 8.10567
R6411 IREF.n1198 IREF.t200 8.10567
R6412 IREF.n1190 IREF.t113 8.10567
R6413 IREF.n124 IREF.t51 8.10567
R6414 IREF.n1260 IREF.t227 8.10567
R6415 IREF.n1266 IREF.t162 8.10567
R6416 IREF.n113 IREF.t154 8.10567
R6417 IREF.n106 IREF.t165 8.10567
R6418 IREF.n101 IREF.t45 8.10567
R6419 IREF.n1287 IREF.t58 8.10567
R6420 IREF.n1196 IREF.t62 8.10567
R6421 IREF.n1195 IREF.t220 8.10567
R6422 IREF.n1245 IREF.t69 8.10567
R6423 IREF.n94 IREF.t198 8.10567
R6424 IREF.n87 IREF.t127 8.10567
R6425 IREF.n45 IREF.t143 8.10567
R6426 IREF.n52 IREF.t169 8.10567
R6427 IREF.n54 IREF.t157 8.10567
R6428 IREF.n58 IREF.t139 8.10567
R6429 IREF.n209 IREF.t156 8.10567
R6430 IREF.n282 IREF.t71 8.10567
R6431 IREF.n276 IREF.t60 8.10567
R6432 IREF.n271 IREF.t208 8.10567
R6433 IREF.n266 IREF.t247 8.10567
R6434 IREF.n326 IREF.t101 8.10567
R6435 IREF.n336 IREF.t174 8.10567
R6436 IREF.n345 IREF.t84 8.10567
R6437 IREF.n354 IREF.t151 8.10567
R6438 IREF.n243 IREF.t218 8.10567
R6439 IREF.n236 IREF.t259 8.10567
R6440 IREF.n231 IREF.t191 8.10567
R6441 IREF.n226 IREF.t236 8.10567
R6442 IREF.n263 IREF.t64 8.10567
R6443 IREF.n262 IREF.t132 8.10567
R6444 IREF.n322 IREF.t122 8.10567
R6445 IREF.n223 IREF.t215 8.10567
R6446 IREF.n216 IREF.t67 8.10567
R6447 IREF.n166 IREF.t110 8.10567
R6448 IREF.n198 IREF.t161 8.10567
R6449 IREF.n189 IREF.t95 8.10567
R6450 IREF.n180 IREF.t225 8.10567
R6451 IREF.n396 IREF.t146 8.10567
R6452 IREF.n531 IREF.t53 8.10567
R6453 IREF.n525 IREF.t263 8.10567
R6454 IREF.n520 IREF.t195 8.10567
R6455 IREF.n549 IREF.t239 8.10567
R6456 IREF.n499 IREF.t94 8.10567
R6457 IREF.n143 IREF.t164 8.10567
R6458 IREF.n145 IREF.t73 8.10567
R6459 IREF.n476 IREF.t136 8.10567
R6460 IREF.n471 IREF.t204 8.10567
R6461 IREF.n155 IREF.t244 8.10567
R6462 IREF.n157 IREF.t175 8.10567
R6463 IREF.n448 IREF.t226 8.10567
R6464 IREF.n513 IREF.t248 8.10567
R6465 IREF.n506 IREF.t105 8.10567
R6466 IREF.n136 IREF.t99 8.10567
R6467 IREF.n444 IREF.t182 8.10567
R6468 IREF.n437 IREF.t252 8.10567
R6469 IREF.n394 IREF.t90 8.10567
R6470 IREF.n400 IREF.t150 8.10567
R6471 IREF.n405 IREF.t86 8.10567
R6472 IREF.n407 IREF.t214 8.10567
R6473 IREF.n591 IREF.t74 8.10567
R6474 IREF.n754 IREF.t196 8.10567
R6475 IREF.n748 IREF.t186 8.10567
R6476 IREF.n743 IREF.t115 8.10567
R6477 IREF.n738 IREF.t163 8.10567
R6478 IREF.n721 IREF.t231 8.10567
R6479 IREF.n710 IREF.t92 8.10567
R6480 IREF.n701 IREF.t212 8.10567
R6481 IREF.n692 IREF.t63 8.10567
R6482 IREF.n576 IREF.t119 8.10567
R6483 IREF.n672 IREF.t171 8.10567
R6484 IREF.n584 IREF.t98 8.10567
R6485 IREF.n588 IREF.t148 8.10567
R6486 IREF.n735 IREF.t190 8.10567
R6487 IREF.n728 IREF.t260 8.10567
R6488 IREF.n560 IREF.t251 8.10567
R6489 IREF.n637 IREF.t117 8.10567
R6490 IREF.n636 IREF.t194 8.10567
R6491 IREF.n647 IREF.t238 8.10567
R6492 IREF.n619 IREF.t78 8.10567
R6493 IREF.n599 IREF.t224 8.10567
R6494 IREF.n603 IREF.t126 8.10567
R6495 IREF.n1161 IREF.t129 8.10567
R6496 IREF.n1155 IREF.t77 8.10567
R6497 IREF.n1148 IREF.t242 8.10567
R6498 IREF.n792 IREF.t180 8.10567
R6499 IREF.n1165 IREF.t257 8.10567
R6500 IREF.n1164 IREF.t199 8.10567
R6501 IREF.n1163 IREF.t262 8.10567
R6502 IREF.n1169 IREF.t103 8.10567
R6503 IREF.n1175 IREF.t209 8.10567
R6504 IREF.n1181 IREF.t221 8.10567
R6505 IREF.n800 IREF.t49 8.10567
R6506 IREF.n802 IREF.t189 8.10567
R6507 IREF.n804 IREF.t178 8.10567
R6508 IREF.n1123 IREF.t177 8.10567
R6509 IREF.n1122 IREF.t112 8.10567
R6510 IREF.n1121 IREF.t120 8.10567
R6511 IREF.n1142 IREF.t172 8.10567
R6512 IREF.n1135 IREF.t183 8.10567
R6513 IREF.n796 IREF.t70 8.10567
R6514 IREF.n798 IREF.t83 8.10567
R6515 IREF.n928 IREF.t91 8.10567
R6516 IREF.n921 IREF.t155 8.10567
R6517 IREF.n915 IREF.t61 8.10567
R6518 IREF.n909 IREF.t128 8.10567
R6519 IREF.n932 IREF.t87 8.10567
R6520 IREF.n931 IREF.t153 8.10567
R6521 IREF.n930 IREF.t147 8.10567
R6522 IREF.n936 IREF.t255 8.10567
R6523 IREF.n935 IREF.t184 8.10567
R6524 IREF.n947 IREF.t232 8.10567
R6525 IREF.n865 IREF.t137 8.10567
R6526 IREF.n874 IREF.t140 8.10567
R6527 IREF.n869 IREF.t82 8.10567
R6528 IREF.n887 IREF.t229 8.10567
R6529 IREF.n886 IREF.t88 8.10567
R6530 IREF.n885 IREF.t125 8.10567
R6531 IREF.n907 IREF.t197 8.10567
R6532 IREF.n900 IREF.t240 8.10567
R6533 IREF.n893 IREF.t170 8.10567
R6534 IREF.n864 IREF.t223 8.10567
R6535 IREF.n851 IREF.t59 8.10567
R6536 IREF.n849 IREF.t124 8.10567
R6537 IREF.n848 IREF.t246 8.10567
R6538 IREF.n992 IREF.t104 8.10567
R6539 IREF.n973 IREF.t75 8.10567
R6540 IREF.n974 IREF.t138 8.10567
R6541 IREF.n975 IREF.t131 8.10567
R6542 IREF.n958 IREF.t230 8.10567
R6543 IREF.n956 IREF.t158 8.10567
R6544 IREF.n955 IREF.t210 8.10567
R6545 IREF.n834 IREF.t109 8.10567
R6546 IREF.n828 IREF.t114 8.10567
R6547 IREF.n822 IREF.t47 8.10567
R6548 IREF.n838 IREF.t222 8.10567
R6549 IREF.n837 IREF.t79 8.10567
R6550 IREF.n836 IREF.t116 8.10567
R6551 IREF.n844 IREF.t167 8.10567
R6552 IREF.n843 IREF.t219 8.10567
R6553 IREF.n1004 IREF.t144 8.10567
R6554 IREF.n1010 IREF.t193 8.10567
R6555 IREF.n1054 IREF.t217 8.10567
R6556 IREF.n1050 IREF.t72 8.10567
R6557 IREF.n1049 IREF.t188 8.10567
R6558 IREF.n1093 IREF.t258 8.10567
R6559 IREF.n1073 IREF.t213 8.10567
R6560 IREF.n1074 IREF.t65 8.10567
R6561 IREF.n1075 IREF.t56 8.10567
R6562 IREF.n1059 IREF.t166 8.10567
R6563 IREF.n1057 IREF.t96 8.10567
R6564 IREF.n1055 IREF.t142 8.10567
R6565 IREF.n1035 IREF.t48 8.10567
R6566 IREF.n1028 IREF.t52 8.10567
R6567 IREF.n1022 IREF.t206 8.10567
R6568 IREF.n1039 IREF.t135 8.10567
R6569 IREF.n1038 IREF.t216 8.10567
R6570 IREF.n1037 IREF.t256 8.10567
R6571 IREF.n1095 IREF.t102 8.10567
R6572 IREF.n1043 IREF.t152 8.10567
R6573 IREF.n1042 IREF.t85 8.10567
R6574 IREF.n1112 IREF.t123 8.10567
R6575 IREF.n1371 IREF.t26 8.10567
R6576 IREF.n1376 IREF.t14 8.10567
R6577 IREF.n1367 IREF.t4 8.10567
R6578 IREF.n1362 IREF.t24 8.10567
R6579 IREF.n1355 IREF.t30 8.10567
R6580 IREF.n1350 IREF.t36 8.10567
R6581 IREF.n21 IREF.t23 6.61324
R6582 IREF.n27 IREF.t9 6.47665
R6583 IREF.n5 IREF.t19 6.43481
R6584 IREF.n19 IREF.t1 6.43476
R6585 IREF.n23 IREF.t11 5.34147
R6586 IREF.n22 IREF.t29 5.34147
R6587 IREF.n182 IREF.n179 4.65575
R6588 IREF.n604 IREF.n602 4.65575
R6589 IREF.n283 IREF.n280 4.64641
R6590 IREF.n755 IREF.n750 4.64641
R6591 IREF.n1143 IREF.n1142 4.64261
R6592 IREF.n994 IREF.n844 4.64261
R6593 IREF.n1363 IREF.n1362 4.64261
R6594 IREF.n59 IREF.n57 4.64
R6595 IREF.n1215 IREF.n1214 4.64
R6596 IREF.n286 IREF.n280 4.64
R6597 IREF.n408 IREF.n406 4.64
R6598 IREF.n533 IREF.n532 4.64
R6599 IREF.n410 IREF.n406 4.64
R6600 IREF.n534 IREF.n533 4.64
R6601 IREF.n756 IREF.n755 4.64
R6602 IREF.n60 IREF.n59 4.64
R6603 IREF.n1216 IREF.n1215 4.64
R6604 IREF.n908 IREF.n907 4.61892
R6605 IREF.n1096 IREF.n1095 4.61892
R6606 IREF.n910 IREF.n909 4.61655
R6607 IREF.n1094 IREF.n1093 4.61655
R6608 IREF.n27 IREF.n26 4.61078
R6609 IREF.n17 IREF.n16 4.61078
R6610 IREF.n13 IREF.n12 4.61078
R6611 IREF.n9 IREF.n8 4.61078
R6612 IREF.n19 IREF.n1 4.61078
R6613 IREF.n35 IREF.n33 4.60951
R6614 IREF.n36 IREF.n35 4.60951
R6615 IREF.n16 IREF.n14 4.60825
R6616 IREF.n12 IREF.n10 4.60825
R6617 IREF.n8 IREF.n5 4.60825
R6618 IREF.n18 IREF.n1 4.60825
R6619 IREF.n1235 IREF.n1196 4.54125
R6620 IREF.n95 IREF.n94 4.54125
R6621 IREF.n514 IREF.n513 4.54125
R6622 IREF.n445 IREF.n444 4.54125
R6623 IREF.n312 IREF.n263 4.53893
R6624 IREF.n224 IREF.n223 4.53893
R6625 IREF.n736 IREF.n735 4.53893
R6626 IREF.n637 IREF.n589 4.53893
R6627 IREF.n310 IREF.n265 4.51011
R6628 IREF.n357 IREF.n356 4.51011
R6629 IREF.n387 IREF.n386 4.51011
R6630 IREF.n782 IREF.n781 4.51011
R6631 IREF.n689 IREF.n574 4.51011
R6632 IREF.n655 IREF.n653 4.51011
R6633 IREF.n325 IREF.n257 4.50691
R6634 IREF.n359 IREF.n358 4.50691
R6635 IREF.n210 IREF.n160 4.50691
R6636 IREF.n722 IREF.n554 4.50691
R6637 IREF.n688 IREF.n687 4.50691
R6638 IREF.n651 IREF.n650 4.50691
R6639 IREF.n34 IREF.n29 4.5005
R6640 IREF.n93 IREF.n42 4.5005
R6641 IREF.n92 IREF.n91 4.5005
R6642 IREF.n90 IREF.n43 4.5005
R6643 IREF.n89 IREF.n88 4.5005
R6644 IREF.n86 IREF.n44 4.5005
R6645 IREF.n85 IREF.n84 4.5005
R6646 IREF.n1237 IREF.n1236 4.5005
R6647 IREF.n1238 IREF.n1194 4.5005
R6648 IREF.n1240 IREF.n1239 4.5005
R6649 IREF.n1241 IREF.n1193 4.5005
R6650 IREF.n1243 IREF.n1242 4.5005
R6651 IREF.n1244 IREF.n1192 4.5005
R6652 IREF.n1270 IREF.n1269 4.5005
R6653 IREF.n114 IREF.n111 4.5005
R6654 IREF.n1274 IREF.n110 4.5005
R6655 IREF.n1275 IREF.n109 4.5005
R6656 IREF.n1276 IREF.n108 4.5005
R6657 IREF.n1279 IREF.n105 4.5005
R6658 IREF.n1280 IREF.n104 4.5005
R6659 IREF.n1281 IREF.n103 4.5005
R6660 IREF.n102 IREF.n99 4.5005
R6661 IREF.n1285 IREF.n98 4.5005
R6662 IREF.n1286 IREF.n97 4.5005
R6663 IREF.n1288 IREF.n96 4.5005
R6664 IREF.n1248 IREF.n1247 4.5005
R6665 IREF.n1191 IREF.n129 4.5005
R6666 IREF.n1252 IREF.n128 4.5005
R6667 IREF.n1253 IREF.n127 4.5005
R6668 IREF.n1254 IREF.n126 4.5005
R6669 IREF.n125 IREF.n122 4.5005
R6670 IREF.n1258 IREF.n121 4.5005
R6671 IREF.n1259 IREF.n120 4.5005
R6672 IREF.n1261 IREF.n119 4.5005
R6673 IREF.n118 IREF.n116 4.5005
R6674 IREF.n1265 IREF.n115 4.5005
R6675 IREF.n1268 IREF.n1267 4.5005
R6676 IREF.n1214 IREF.n1212 4.5005
R6677 IREF.n1218 IREF.n1211 4.5005
R6678 IREF.n1219 IREF.n1210 4.5005
R6679 IREF.n1220 IREF.n1209 4.5005
R6680 IREF.n1223 IREF.n1206 4.5005
R6681 IREF.n1224 IREF.n1205 4.5005
R6682 IREF.n1225 IREF.n1204 4.5005
R6683 IREF.n1228 IREF.n1201 4.5005
R6684 IREF.n1229 IREF.n1200 4.5005
R6685 IREF.n1230 IREF.n1197 4.5005
R6686 IREF.n1234 IREF.n1233 4.5005
R6687 IREF.n82 IREF.n81 4.5005
R6688 IREF.n79 IREF.n46 4.5005
R6689 IREF.n73 IREF.n47 4.5005
R6690 IREF.n75 IREF.n74 4.5005
R6691 IREF.n72 IREF.n49 4.5005
R6692 IREF.n71 IREF.n70 4.5005
R6693 IREF.n51 IREF.n50 4.5005
R6694 IREF.n66 IREF.n65 4.5005
R6695 IREF.n64 IREF.n63 4.5005
R6696 IREF.n62 IREF.n55 4.5005
R6697 IREF.n57 IREF.n56 4.5005
R6698 IREF.n222 IREF.n163 4.5005
R6699 IREF.n221 IREF.n220 4.5005
R6700 IREF.n219 IREF.n164 4.5005
R6701 IREF.n218 IREF.n217 4.5005
R6702 IREF.n215 IREF.n165 4.5005
R6703 IREF.n214 IREF.n213 4.5005
R6704 IREF.n314 IREF.n313 4.5005
R6705 IREF.n315 IREF.n261 4.5005
R6706 IREF.n317 IREF.n316 4.5005
R6707 IREF.n318 IREF.n260 4.5005
R6708 IREF.n320 IREF.n319 4.5005
R6709 IREF.n321 IREF.n259 4.5005
R6710 IREF.n386 IREF.n385 4.5005
R6711 IREF.n384 IREF.n383 4.5005
R6712 IREF.n227 IREF.n225 4.5005
R6713 IREF.n378 IREF.n377 4.5005
R6714 IREF.n376 IREF.n375 4.5005
R6715 IREF.n232 IREF.n230 4.5005
R6716 IREF.n370 IREF.n369 4.5005
R6717 IREF.n368 IREF.n367 4.5005
R6718 IREF.n237 IREF.n235 4.5005
R6719 IREF.n241 IREF.n239 4.5005
R6720 IREF.n362 IREF.n361 4.5005
R6721 IREF.n360 IREF.n359 4.5005
R6722 IREF.n356 IREF.n242 4.5005
R6723 IREF.n353 IREF.n352 4.5005
R6724 IREF.n351 IREF.n350 4.5005
R6725 IREF.n247 IREF.n246 4.5005
R6726 IREF.n344 IREF.n343 4.5005
R6727 IREF.n342 IREF.n341 4.5005
R6728 IREF.n252 IREF.n251 4.5005
R6729 IREF.n335 IREF.n334 4.5005
R6730 IREF.n333 IREF.n332 4.5005
R6731 IREF.n331 IREF.n255 4.5005
R6732 IREF.n258 IREF.n256 4.5005
R6733 IREF.n325 IREF.n324 4.5005
R6734 IREF.n311 IREF.n310 4.5005
R6735 IREF.n268 IREF.n264 4.5005
R6736 IREF.n305 IREF.n304 4.5005
R6737 IREF.n303 IREF.n302 4.5005
R6738 IREF.n273 IREF.n270 4.5005
R6739 IREF.n297 IREF.n296 4.5005
R6740 IREF.n295 IREF.n294 4.5005
R6741 IREF.n278 IREF.n275 4.5005
R6742 IREF.n289 IREF.n288 4.5005
R6743 IREF.n287 IREF.n279 4.5005
R6744 IREF.n286 IREF.n285 4.5005
R6745 IREF.n182 IREF.n181 4.5005
R6746 IREF.n184 IREF.n183 4.5005
R6747 IREF.n176 IREF.n175 4.5005
R6748 IREF.n191 IREF.n190 4.5005
R6749 IREF.n193 IREF.n192 4.5005
R6750 IREF.n172 IREF.n171 4.5005
R6751 IREF.n201 IREF.n200 4.5005
R6752 IREF.n202 IREF.n170 4.5005
R6753 IREF.n204 IREF.n203 4.5005
R6754 IREF.n168 IREF.n167 4.5005
R6755 IREF.n211 IREF.n210 4.5005
R6756 IREF.n178 IREF.n177 4.5005
R6757 IREF.n186 IREF.n185 4.5005
R6758 IREF.n188 IREF.n187 4.5005
R6759 IREF.n174 IREF.n173 4.5005
R6760 IREF.n195 IREF.n194 4.5005
R6761 IREF.n197 IREF.n196 4.5005
R6762 IREF.n199 IREF.n169 4.5005
R6763 IREF.n206 IREF.n205 4.5005
R6764 IREF.n208 IREF.n207 4.5005
R6765 IREF.n162 IREF.n161 4.5005
R6766 IREF.n382 IREF.n381 4.5005
R6767 IREF.n380 IREF.n379 4.5005
R6768 IREF.n229 IREF.n228 4.5005
R6769 IREF.n374 IREF.n373 4.5005
R6770 IREF.n372 IREF.n371 4.5005
R6771 IREF.n234 IREF.n233 4.5005
R6772 IREF.n366 IREF.n365 4.5005
R6773 IREF.n364 IREF.n363 4.5005
R6774 IREF.n240 IREF.n238 4.5005
R6775 IREF.n355 IREF.n244 4.5005
R6776 IREF.n248 IREF.n245 4.5005
R6777 IREF.n349 IREF.n348 4.5005
R6778 IREF.n347 IREF.n346 4.5005
R6779 IREF.n250 IREF.n249 4.5005
R6780 IREF.n340 IREF.n339 4.5005
R6781 IREF.n338 IREF.n337 4.5005
R6782 IREF.n254 IREF.n253 4.5005
R6783 IREF.n330 IREF.n329 4.5005
R6784 IREF.n328 IREF.n327 4.5005
R6785 IREF.n309 IREF.n308 4.5005
R6786 IREF.n307 IREF.n306 4.5005
R6787 IREF.n269 IREF.n267 4.5005
R6788 IREF.n301 IREF.n300 4.5005
R6789 IREF.n299 IREF.n298 4.5005
R6790 IREF.n274 IREF.n272 4.5005
R6791 IREF.n293 IREF.n292 4.5005
R6792 IREF.n291 IREF.n290 4.5005
R6793 IREF.n281 IREF.n277 4.5005
R6794 IREF.n284 IREF.n283 4.5005
R6795 IREF.n443 IREF.n391 4.5005
R6796 IREF.n442 IREF.n441 4.5005
R6797 IREF.n440 IREF.n392 4.5005
R6798 IREF.n439 IREF.n438 4.5005
R6799 IREF.n436 IREF.n393 4.5005
R6800 IREF.n435 IREF.n434 4.5005
R6801 IREF.n512 IREF.n133 4.5005
R6802 IREF.n511 IREF.n510 4.5005
R6803 IREF.n509 IREF.n134 4.5005
R6804 IREF.n508 IREF.n507 4.5005
R6805 IREF.n505 IREF.n135 4.5005
R6806 IREF.n504 IREF.n503 4.5005
R6807 IREF.n473 IREF.n472 4.5005
R6808 IREF.n470 IREF.n149 4.5005
R6809 IREF.n464 IREF.n150 4.5005
R6810 IREF.n466 IREF.n465 4.5005
R6811 IREF.n463 IREF.n152 4.5005
R6812 IREF.n462 IREF.n461 4.5005
R6813 IREF.n154 IREF.n153 4.5005
R6814 IREF.n457 IREF.n456 4.5005
R6815 IREF.n455 IREF.n454 4.5005
R6816 IREF.n453 IREF.n158 4.5005
R6817 IREF.n446 IREF.n159 4.5005
R6818 IREF.n449 IREF.n447 4.5005
R6819 IREF.n501 IREF.n500 4.5005
R6820 IREF.n498 IREF.n137 4.5005
R6821 IREF.n492 IREF.n138 4.5005
R6822 IREF.n494 IREF.n493 4.5005
R6823 IREF.n491 IREF.n140 4.5005
R6824 IREF.n490 IREF.n489 4.5005
R6825 IREF.n142 IREF.n141 4.5005
R6826 IREF.n485 IREF.n484 4.5005
R6827 IREF.n483 IREF.n482 4.5005
R6828 IREF.n481 IREF.n146 4.5005
R6829 IREF.n474 IREF.n147 4.5005
R6830 IREF.n477 IREF.n475 4.5005
R6831 IREF.n532 IREF.n530 4.5005
R6832 IREF.n536 IREF.n529 4.5005
R6833 IREF.n537 IREF.n528 4.5005
R6834 IREF.n538 IREF.n527 4.5005
R6835 IREF.n541 IREF.n524 4.5005
R6836 IREF.n542 IREF.n523 4.5005
R6837 IREF.n543 IREF.n522 4.5005
R6838 IREF.n521 IREF.n518 4.5005
R6839 IREF.n547 IREF.n517 4.5005
R6840 IREF.n548 IREF.n516 4.5005
R6841 IREF.n550 IREF.n515 4.5005
R6842 IREF.n432 IREF.n431 4.5005
R6843 IREF.n428 IREF.n395 4.5005
R6844 IREF.n427 IREF.n426 4.5005
R6845 IREF.n425 IREF.n398 4.5005
R6846 IREF.n424 IREF.n423 4.5005
R6847 IREF.n419 IREF.n399 4.5005
R6848 IREF.n418 IREF.n417 4.5005
R6849 IREF.n416 IREF.n402 4.5005
R6850 IREF.n415 IREF.n414 4.5005
R6851 IREF.n404 IREF.n403 4.5005
R6852 IREF.n409 IREF.n408 4.5005
R6853 IREF.n410 IREF.n409 4.5005
R6854 IREF.n411 IREF.n404 4.5005
R6855 IREF.n414 IREF.n413 4.5005
R6856 IREF.n412 IREF.n402 4.5005
R6857 IREF.n418 IREF.n401 4.5005
R6858 IREF.n420 IREF.n419 4.5005
R6859 IREF.n423 IREF.n422 4.5005
R6860 IREF.n421 IREF.n398 4.5005
R6861 IREF.n427 IREF.n397 4.5005
R6862 IREF.n429 IREF.n428 4.5005
R6863 IREF.n431 IREF.n430 4.5005
R6864 IREF.n450 IREF.n449 4.5005
R6865 IREF.n451 IREF.n159 4.5005
R6866 IREF.n453 IREF.n452 4.5005
R6867 IREF.n454 IREF.n156 4.5005
R6868 IREF.n458 IREF.n457 4.5005
R6869 IREF.n459 IREF.n154 4.5005
R6870 IREF.n461 IREF.n460 4.5005
R6871 IREF.n152 IREF.n151 4.5005
R6872 IREF.n467 IREF.n466 4.5005
R6873 IREF.n468 IREF.n150 4.5005
R6874 IREF.n470 IREF.n469 4.5005
R6875 IREF.n472 IREF.n148 4.5005
R6876 IREF.n478 IREF.n477 4.5005
R6877 IREF.n479 IREF.n147 4.5005
R6878 IREF.n481 IREF.n480 4.5005
R6879 IREF.n482 IREF.n144 4.5005
R6880 IREF.n486 IREF.n485 4.5005
R6881 IREF.n487 IREF.n142 4.5005
R6882 IREF.n489 IREF.n488 4.5005
R6883 IREF.n140 IREF.n139 4.5005
R6884 IREF.n495 IREF.n494 4.5005
R6885 IREF.n496 IREF.n138 4.5005
R6886 IREF.n498 IREF.n497 4.5005
R6887 IREF.n500 IREF.n131 4.5005
R6888 IREF.n551 IREF.n550 4.5005
R6889 IREF.n548 IREF.n132 4.5005
R6890 IREF.n547 IREF.n546 4.5005
R6891 IREF.n545 IREF.n518 4.5005
R6892 IREF.n544 IREF.n543 4.5005
R6893 IREF.n542 IREF.n519 4.5005
R6894 IREF.n541 IREF.n540 4.5005
R6895 IREF.n539 IREF.n538 4.5005
R6896 IREF.n537 IREF.n526 4.5005
R6897 IREF.n536 IREF.n535 4.5005
R6898 IREF.n534 IREF.n530 4.5005
R6899 IREF.n639 IREF.n638 4.5005
R6900 IREF.n640 IREF.n635 4.5005
R6901 IREF.n642 IREF.n641 4.5005
R6902 IREF.n643 IREF.n634 4.5005
R6903 IREF.n645 IREF.n644 4.5005
R6904 IREF.n646 IREF.n633 4.5005
R6905 IREF.n734 IREF.n557 4.5005
R6906 IREF.n733 IREF.n732 4.5005
R6907 IREF.n731 IREF.n558 4.5005
R6908 IREF.n730 IREF.n729 4.5005
R6909 IREF.n727 IREF.n559 4.5005
R6910 IREF.n726 IREF.n725 4.5005
R6911 IREF.n656 IREF.n655 4.5005
R6912 IREF.n658 IREF.n657 4.5005
R6913 IREF.n586 IREF.n585 4.5005
R6914 IREF.n665 IREF.n664 4.5005
R6915 IREF.n667 IREF.n666 4.5005
R6916 IREF.n582 IREF.n581 4.5005
R6917 IREF.n675 IREF.n674 4.5005
R6918 IREF.n676 IREF.n580 4.5005
R6919 IREF.n678 IREF.n677 4.5005
R6920 IREF.n578 IREF.n577 4.5005
R6921 IREF.n685 IREF.n684 4.5005
R6922 IREF.n687 IREF.n686 4.5005
R6923 IREF.n574 IREF.n573 4.5005
R6924 IREF.n694 IREF.n693 4.5005
R6925 IREF.n696 IREF.n695 4.5005
R6926 IREF.n570 IREF.n569 4.5005
R6927 IREF.n703 IREF.n702 4.5005
R6928 IREF.n705 IREF.n704 4.5005
R6929 IREF.n566 IREF.n565 4.5005
R6930 IREF.n713 IREF.n712 4.5005
R6931 IREF.n714 IREF.n564 4.5005
R6932 IREF.n716 IREF.n715 4.5005
R6933 IREF.n562 IREF.n561 4.5005
R6934 IREF.n723 IREF.n722 4.5005
R6935 IREF.n781 IREF.n780 4.5005
R6936 IREF.n779 IREF.n778 4.5005
R6937 IREF.n739 IREF.n737 4.5005
R6938 IREF.n773 IREF.n772 4.5005
R6939 IREF.n771 IREF.n770 4.5005
R6940 IREF.n744 IREF.n742 4.5005
R6941 IREF.n765 IREF.n764 4.5005
R6942 IREF.n763 IREF.n762 4.5005
R6943 IREF.n749 IREF.n747 4.5005
R6944 IREF.n753 IREF.n751 4.5005
R6945 IREF.n757 IREF.n756 4.5005
R6946 IREF.n605 IREF.n604 4.5005
R6947 IREF.n601 IREF.n600 4.5005
R6948 IREF.n612 IREF.n611 4.5005
R6949 IREF.n614 IREF.n613 4.5005
R6950 IREF.n597 IREF.n596 4.5005
R6951 IREF.n622 IREF.n621 4.5005
R6952 IREF.n623 IREF.n595 4.5005
R6953 IREF.n625 IREF.n624 4.5005
R6954 IREF.n593 IREF.n592 4.5005
R6955 IREF.n632 IREF.n631 4.5005
R6956 IREF.n650 IREF.n649 4.5005
R6957 IREF.n607 IREF.n606 4.5005
R6958 IREF.n609 IREF.n608 4.5005
R6959 IREF.n610 IREF.n598 4.5005
R6960 IREF.n616 IREF.n615 4.5005
R6961 IREF.n618 IREF.n617 4.5005
R6962 IREF.n620 IREF.n594 4.5005
R6963 IREF.n627 IREF.n626 4.5005
R6964 IREF.n629 IREF.n628 4.5005
R6965 IREF.n630 IREF.n590 4.5005
R6966 IREF.n654 IREF.n587 4.5005
R6967 IREF.n660 IREF.n659 4.5005
R6968 IREF.n662 IREF.n661 4.5005
R6969 IREF.n663 IREF.n583 4.5005
R6970 IREF.n669 IREF.n668 4.5005
R6971 IREF.n671 IREF.n670 4.5005
R6972 IREF.n673 IREF.n579 4.5005
R6973 IREF.n680 IREF.n679 4.5005
R6974 IREF.n682 IREF.n681 4.5005
R6975 IREF.n683 IREF.n575 4.5005
R6976 IREF.n691 IREF.n690 4.5005
R6977 IREF.n572 IREF.n571 4.5005
R6978 IREF.n698 IREF.n697 4.5005
R6979 IREF.n700 IREF.n699 4.5005
R6980 IREF.n568 IREF.n567 4.5005
R6981 IREF.n707 IREF.n706 4.5005
R6982 IREF.n709 IREF.n708 4.5005
R6983 IREF.n711 IREF.n563 4.5005
R6984 IREF.n718 IREF.n717 4.5005
R6985 IREF.n720 IREF.n719 4.5005
R6986 IREF.n556 IREF.n555 4.5005
R6987 IREF.n777 IREF.n776 4.5005
R6988 IREF.n775 IREF.n774 4.5005
R6989 IREF.n741 IREF.n740 4.5005
R6990 IREF.n769 IREF.n768 4.5005
R6991 IREF.n767 IREF.n766 4.5005
R6992 IREF.n746 IREF.n745 4.5005
R6993 IREF.n761 IREF.n760 4.5005
R6994 IREF.n759 IREF.n758 4.5005
R6995 IREF.n752 IREF.n750 4.5005
R6996 IREF.n60 IREF.n56 4.5005
R6997 IREF.n62 IREF.n61 4.5005
R6998 IREF.n63 IREF.n53 4.5005
R6999 IREF.n67 IREF.n66 4.5005
R7000 IREF.n68 IREF.n51 4.5005
R7001 IREF.n70 IREF.n69 4.5005
R7002 IREF.n49 IREF.n48 4.5005
R7003 IREF.n76 IREF.n75 4.5005
R7004 IREF.n77 IREF.n47 4.5005
R7005 IREF.n79 IREF.n78 4.5005
R7006 IREF.n81 IREF.n40 4.5005
R7007 IREF.n1289 IREF.n1288 4.5005
R7008 IREF.n1286 IREF.n41 4.5005
R7009 IREF.n1285 IREF.n1284 4.5005
R7010 IREF.n1283 IREF.n99 4.5005
R7011 IREF.n1282 IREF.n1281 4.5005
R7012 IREF.n1280 IREF.n100 4.5005
R7013 IREF.n1279 IREF.n1278 4.5005
R7014 IREF.n1277 IREF.n1276 4.5005
R7015 IREF.n1275 IREF.n107 4.5005
R7016 IREF.n1274 IREF.n1273 4.5005
R7017 IREF.n1272 IREF.n111 4.5005
R7018 IREF.n1271 IREF.n1270 4.5005
R7019 IREF.n1267 IREF.n112 4.5005
R7020 IREF.n1265 IREF.n1264 4.5005
R7021 IREF.n1263 IREF.n116 4.5005
R7022 IREF.n1262 IREF.n1261 4.5005
R7023 IREF.n1259 IREF.n117 4.5005
R7024 IREF.n1258 IREF.n1257 4.5005
R7025 IREF.n1256 IREF.n122 4.5005
R7026 IREF.n1255 IREF.n1254 4.5005
R7027 IREF.n1253 IREF.n123 4.5005
R7028 IREF.n1252 IREF.n1251 4.5005
R7029 IREF.n1250 IREF.n129 4.5005
R7030 IREF.n1249 IREF.n1248 4.5005
R7031 IREF.n1233 IREF.n1232 4.5005
R7032 IREF.n1231 IREF.n1230 4.5005
R7033 IREF.n1229 IREF.n1199 4.5005
R7034 IREF.n1228 IREF.n1227 4.5005
R7035 IREF.n1226 IREF.n1225 4.5005
R7036 IREF.n1224 IREF.n1203 4.5005
R7037 IREF.n1223 IREF.n1222 4.5005
R7038 IREF.n1221 IREF.n1220 4.5005
R7039 IREF.n1219 IREF.n1208 4.5005
R7040 IREF.n1218 IREF.n1217 4.5005
R7041 IREF.n1216 IREF.n1212 4.5005
R7042 IREF.n872 IREF.n871 4.5005
R7043 IREF.n873 IREF.n868 4.5005
R7044 IREF.n876 IREF.n875 4.5005
R7045 IREF.n877 IREF.n867 4.5005
R7046 IREF.n879 IREF.n878 4.5005
R7047 IREF.n880 IREF.n866 4.5005
R7048 IREF.n882 IREF.n881 4.5005
R7049 IREF.n884 IREF.n883 4.5005
R7050 IREF.n889 IREF.n888 4.5005
R7051 IREF.n891 IREF.n890 4.5005
R7052 IREF.n892 IREF.n863 4.5005
R7053 IREF.n895 IREF.n894 4.5005
R7054 IREF.n896 IREF.n862 4.5005
R7055 IREF.n898 IREF.n897 4.5005
R7056 IREF.n899 IREF.n861 4.5005
R7057 IREF.n902 IREF.n901 4.5005
R7058 IREF.n903 IREF.n860 4.5005
R7059 IREF.n905 IREF.n904 4.5005
R7060 IREF.n906 IREF.n859 4.5005
R7061 IREF.n911 IREF.n858 4.5005
R7062 IREF.n913 IREF.n912 4.5005
R7063 IREF.n914 IREF.n857 4.5005
R7064 IREF.n917 IREF.n916 4.5005
R7065 IREF.n918 IREF.n856 4.5005
R7066 IREF.n920 IREF.n919 4.5005
R7067 IREF.n922 IREF.n855 4.5005
R7068 IREF.n924 IREF.n923 4.5005
R7069 IREF.n925 IREF.n854 4.5005
R7070 IREF.n927 IREF.n926 4.5005
R7071 IREF.n929 IREF.n852 4.5005
R7072 IREF.n949 IREF.n948 4.5005
R7073 IREF.n946 IREF.n853 4.5005
R7074 IREF.n945 IREF.n944 4.5005
R7075 IREF.n943 IREF.n933 4.5005
R7076 IREF.n942 IREF.n941 4.5005
R7077 IREF.n940 IREF.n934 4.5005
R7078 IREF.n939 IREF.n938 4.5005
R7079 IREF.n835 IREF.n817 4.5005
R7080 IREF.n833 IREF.n832 4.5005
R7081 IREF.n831 IREF.n819 4.5005
R7082 IREF.n830 IREF.n829 4.5005
R7083 IREF.n827 IREF.n820 4.5005
R7084 IREF.n826 IREF.n825 4.5005
R7085 IREF.n824 IREF.n821 4.5005
R7086 IREF.n1013 IREF.n1012 4.5005
R7087 IREF.n1011 IREF.n818 4.5005
R7088 IREF.n1009 IREF.n1008 4.5005
R7089 IREF.n1007 IREF.n839 4.5005
R7090 IREF.n1006 IREF.n1005 4.5005
R7091 IREF.n1003 IREF.n840 4.5005
R7092 IREF.n1002 IREF.n1001 4.5005
R7093 IREF.n1000 IREF.n841 4.5005
R7094 IREF.n999 IREF.n998 4.5005
R7095 IREF.n997 IREF.n842 4.5005
R7096 IREF.n996 IREF.n995 4.5005
R7097 IREF.n977 IREF.n976 4.5005
R7098 IREF.n979 IREF.n978 4.5005
R7099 IREF.n980 IREF.n850 4.5005
R7100 IREF.n982 IREF.n981 4.5005
R7101 IREF.n984 IREF.n983 4.5005
R7102 IREF.n985 IREF.n847 4.5005
R7103 IREF.n987 IREF.n986 4.5005
R7104 IREF.n988 IREF.n846 4.5005
R7105 IREF.n990 IREF.n989 4.5005
R7106 IREF.n991 IREF.n845 4.5005
R7107 IREF.n972 IREF.n971 4.5005
R7108 IREF.n970 IREF.n953 4.5005
R7109 IREF.n969 IREF.n968 4.5005
R7110 IREF.n967 IREF.n954 4.5005
R7111 IREF.n966 IREF.n965 4.5005
R7112 IREF.n964 IREF.n963 4.5005
R7113 IREF.n962 IREF.n957 4.5005
R7114 IREF.n961 IREF.n960 4.5005
R7115 IREF.n1024 IREF.n1023 4.5005
R7116 IREF.n1025 IREF.n1020 4.5005
R7117 IREF.n1027 IREF.n1026 4.5005
R7118 IREF.n1029 IREF.n1019 4.5005
R7119 IREF.n1031 IREF.n1030 4.5005
R7120 IREF.n1032 IREF.n1018 4.5005
R7121 IREF.n1034 IREF.n1033 4.5005
R7122 IREF.n1036 IREF.n1016 4.5005
R7123 IREF.n1114 IREF.n1113 4.5005
R7124 IREF.n1111 IREF.n1017 4.5005
R7125 IREF.n1110 IREF.n1109 4.5005
R7126 IREF.n1108 IREF.n1040 4.5005
R7127 IREF.n1107 IREF.n1106 4.5005
R7128 IREF.n1105 IREF.n1041 4.5005
R7129 IREF.n1104 IREF.n1103 4.5005
R7130 IREF.n1102 IREF.n1101 4.5005
R7131 IREF.n1100 IREF.n1044 4.5005
R7132 IREF.n1099 IREF.n1098 4.5005
R7133 IREF.n1097 IREF.n1045 4.5005
R7134 IREF.n1092 IREF.n1046 4.5005
R7135 IREF.n1091 IREF.n1090 4.5005
R7136 IREF.n1089 IREF.n1047 4.5005
R7137 IREF.n1088 IREF.n1087 4.5005
R7138 IREF.n1086 IREF.n1048 4.5005
R7139 IREF.n1085 IREF.n1084 4.5005
R7140 IREF.n1083 IREF.n1082 4.5005
R7141 IREF.n1081 IREF.n1051 4.5005
R7142 IREF.n1080 IREF.n1079 4.5005
R7143 IREF.n1078 IREF.n1052 4.5005
R7144 IREF.n1077 IREF.n1076 4.5005
R7145 IREF.n1072 IREF.n1071 4.5005
R7146 IREF.n1070 IREF.n1069 4.5005
R7147 IREF.n1068 IREF.n1056 4.5005
R7148 IREF.n1067 IREF.n1066 4.5005
R7149 IREF.n1065 IREF.n1064 4.5005
R7150 IREF.n1063 IREF.n1058 4.5005
R7151 IREF.n1062 IREF.n1061 4.5005
R7152 IREF.n1120 IREF.n1119 4.5005
R7153 IREF.n815 IREF.n814 4.5005
R7154 IREF.n813 IREF.n801 4.5005
R7155 IREF.n812 IREF.n811 4.5005
R7156 IREF.n810 IREF.n809 4.5005
R7157 IREF.n808 IREF.n803 4.5005
R7158 IREF.n807 IREF.n806 4.5005
R7159 IREF.n1124 IREF.n799 4.5005
R7160 IREF.n1126 IREF.n1125 4.5005
R7161 IREF.n1128 IREF.n1127 4.5005
R7162 IREF.n1129 IREF.n797 4.5005
R7163 IREF.n1131 IREF.n1130 4.5005
R7164 IREF.n1133 IREF.n1132 4.5005
R7165 IREF.n1134 IREF.n795 4.5005
R7166 IREF.n1137 IREF.n1136 4.5005
R7167 IREF.n1138 IREF.n794 4.5005
R7168 IREF.n1140 IREF.n1139 4.5005
R7169 IREF.n1141 IREF.n793 4.5005
R7170 IREF.n1162 IREF.n786 4.5005
R7171 IREF.n1160 IREF.n1159 4.5005
R7172 IREF.n1158 IREF.n788 4.5005
R7173 IREF.n1157 IREF.n1156 4.5005
R7174 IREF.n1154 IREF.n789 4.5005
R7175 IREF.n1153 IREF.n1152 4.5005
R7176 IREF.n1151 IREF.n790 4.5005
R7177 IREF.n1150 IREF.n1149 4.5005
R7178 IREF.n1147 IREF.n791 4.5005
R7179 IREF.n1146 IREF.n1145 4.5005
R7180 IREF.n1184 IREF.n1183 4.5005
R7181 IREF.n1182 IREF.n787 4.5005
R7182 IREF.n1180 IREF.n1179 4.5005
R7183 IREF.n1178 IREF.n1166 4.5005
R7184 IREF.n1177 IREF.n1176 4.5005
R7185 IREF.n1174 IREF.n1167 4.5005
R7186 IREF.n1173 IREF.n1172 4.5005
R7187 IREF.n1171 IREF.n1168 4.5005
R7188 IREF.n1353 IREF.n1352 4.5005
R7189 IREF.n1354 IREF.n1349 4.5005
R7190 IREF.n1357 IREF.n1356 4.5005
R7191 IREF.n1358 IREF.n1348 4.5005
R7192 IREF.n1360 IREF.n1359 4.5005
R7193 IREF.n1361 IREF.n1347 4.5005
R7194 IREF.n1379 IREF.n1378 4.5005
R7195 IREF.n1377 IREF.n1368 4.5005
R7196 IREF.n1376 IREF.n1375 4.5005
R7197 IREF.n1374 IREF.n1369 4.5005
R7198 IREF.n1373 IREF.n1372 4.5005
R7199 IREF.n7 IREF.n4 4.5005
R7200 IREF.n11 IREF.n3 4.5005
R7201 IREF.n15 IREF.n2 4.5005
R7202 IREF.n1387 IREF.n1386 4.5005
R7203 IREF.n1187 IREF.n38 3.97759
R7204 IREF.n21 IREF.n20 3.87147
R7205 IREF.n34 IREF.t35 3.86699
R7206 IREF.n15 IREF.t5 3.83383
R7207 IREF.n11 IREF.t25 3.83383
R7208 IREF.n35 IREF.t7 3.66094
R7209 IREF.n994 IREF.n993 3.03856
R7210 IREF.n1144 IREF.n1143 3.03856
R7211 IREF.n1269 IREF.n1268 3.0245
R7212 IREF.n360 IREF.n242 3.0245
R7213 IREF.n475 IREF.n473 3.0245
R7214 IREF.n478 IREF.n148 3.0245
R7215 IREF.n686 IREF.n573 3.0245
R7216 IREF.n1271 IREF.n112 3.0245
R7217 IREF.n910 IREF.n908 3.0245
R7218 IREF.n1096 IREF.n1094 3.0245
R7219 IREF.n358 IREF.n357 2.96825
R7220 IREF.n689 IREF.n688 2.96825
R7221 IREF.n37 IREF.n36 2.94838
R7222 IREF.n33 IREF.n32 2.60059
R7223 IREF.n23 IREF.n22 2.51878
R7224 IREF.n37 IREF.n28 2.44398
R7225 IREF.n179 IREF.n177 2.41967
R7226 IREF.n607 IREF.n602 2.41967
R7227 IREF.n26 IREF.n25 2.40646
R7228 IREF.n32 IREF.n30 2.39895
R7229 IREF.n7 IREF.n6 2.36383
R7230 IREF.n1015 IREF.n816 2.30989
R7231 IREF.n951 IREF.n950 2.30989
R7232 IREF IREF.n0 2.28212
R7233 IREF.n1144 IREF.n792 2.25752
R7234 IREF.n993 IREF.n992 2.25752
R7235 IREF.n1380 IREF.n1367 2.25278
R7236 IREF.n14 IREF.n13 2.246
R7237 IREF.n26 IREF.n24 2.24358
R7238 IREF.n1246 IREF.n1245 2.22849
R7239 IREF.n83 IREF.n45 2.22849
R7240 IREF.n502 IREF.n136 2.22849
R7241 IREF.n433 IREF.n394 2.22849
R7242 IREF.n323 IREF.n322 2.22782
R7243 IREF.n212 IREF.n166 2.22782
R7244 IREF.n724 IREF.n560 2.22782
R7245 IREF.n648 IREF.n647 2.22782
R7246 IREF.n32 IREF.n31 2.19216
R7247 IREF.n883 IREF.n816 2.18975
R7248 IREF.n950 IREF.n852 2.18975
R7249 IREF.n1115 IREF.n1016 2.18975
R7250 IREF.n1077 IREF.n1053 2.18975
R7251 IREF.n1014 IREF.n817 2.16725
R7252 IREF.n977 IREF.n952 2.16725
R7253 IREF.n1119 IREF.n1118 2.16725
R7254 IREF.n1185 IREF.n786 2.16725
R7255 IREF.n450 IREF.n390 2.102
R7256 IREF.n552 IREF.n551 2.102
R7257 IREF.n1290 IREF.n1289 2.102
R7258 IREF.n1232 IREF.n1189 2.102
R7259 IREF.n389 IREF.n388 2.07182
R7260 IREF.n553 IREF.n130 2.07182
R7261 IREF.n388 IREF.n387 2.06825
R7262 IREF.n265 IREF.n130 2.06825
R7263 IREF.n653 IREF.n652 2.06825
R7264 IREF.n783 IREF.n782 2.06825
R7265 IREF.n1187 IREF.n1186 2.01366
R7266 IREF.n1384 IREF.n1383 1.91821
R7267 IREF.n1313 IREF.n1302 1.61908
R7268 IREF.n1292 IREF.n1291 1.53101
R7269 IREF.n1188 IREF.n1187 1.53101
R7270 IREF.n652 IREF.n39 1.5005
R7271 IREF.n390 IREF.n389 1.5005
R7272 IREF.n1291 IREF.n1290 1.5005
R7273 IREF.n1189 IREF.n1188 1.5005
R7274 IREF.n784 IREF.n783 1.5005
R7275 IREF.n553 IREF.n552 1.5005
R7276 IREF.n1116 IREF.n1115 1.5005
R7277 IREF.n1015 IREF.n1014 1.5005
R7278 IREF.n1118 IREF.n1117 1.5005
R7279 IREF.n1186 IREF.n1185 1.5005
R7280 IREF.n1053 IREF.n785 1.5005
R7281 IREF.n952 IREF.n951 1.5005
R7282 IREF.n1346 IREF.n1345 1.5005
R7283 IREF.n1335 IREF.n1334 1.5005
R7284 IREF.n1382 IREF.n1381 1.5005
R7285 IREF.n1324 IREF.n1323 1.5005
R7286 IREF.n1313 IREF.n1312 1.5005
R7287 IREF.n1385 IREF.n1384 1.5005
R7288 IREF.n389 IREF.n39 1.47516
R7289 IREF.n784 IREF.n553 1.47516
R7290 IREF.n0 IREF.t15 1.4705
R7291 IREF.n0 IREF.t27 1.4705
R7292 IREF.n25 IREF.t21 1.4705
R7293 IREF.n25 IREF.t33 1.4705
R7294 IREF.n20 IREF.t43 1.4705
R7295 IREF.n20 IREF.t41 1.4705
R7296 IREF.n30 IREF.t3 1.4705
R7297 IREF.n30 IREF.t39 1.4705
R7298 IREF.n31 IREF.t17 1.4705
R7299 IREF.n31 IREF.t13 1.4705
R7300 IREF.n6 IREF.t37 1.4705
R7301 IREF.n6 IREF.t31 1.4705
R7302 IREF.n1383 IREF.n1382 1.42915
R7303 IREF.n1117 IREF.n38 1.41182
R7304 IREF.n960 IREF.n959 1.392
R7305 IREF.n1171 IREF.n1170 1.392
R7306 IREF.n871 IREF.n870 1.38741
R7307 IREF.n1024 IREF.n1021 1.38741
R7308 IREF.n22 IREF.n21 1.27228
R7309 IREF.n948 IREF.n932 1.24866
R7310 IREF.n888 IREF.n887 1.24866
R7311 IREF.n1073 IREF.n1072 1.24866
R7312 IREF.n1113 IREF.n1039 1.24866
R7313 IREF.n930 IREF.n929 1.24629
R7314 IREF.n885 IREF.n884 1.24629
R7315 IREF.n1076 IREF.n1075 1.24629
R7316 IREF.n1037 IREF.n1036 1.24629
R7317 IREF.n1116 IREF.n1015 1.23709
R7318 IREF.n951 IREF.n785 1.23709
R7319 IREF.n1163 IREF.n1162 1.22261
R7320 IREF.n1121 IREF.n1120 1.22261
R7321 IREF.n976 IREF.n975 1.22261
R7322 IREF.n836 IREF.n835 1.22261
R7323 IREF.n1183 IREF.n1165 1.21313
R7324 IREF.n1124 IREF.n1123 1.21313
R7325 IREF.n973 IREF.n972 1.21313
R7326 IREF.n1012 IREF.n838 1.21313
R7327 IREF.n24 IREF.n23 1.20609
R7328 IREF.n824 IREF.n823 1.12904
R7329 IREF.n806 IREF.n805 1.12904
R7330 IREF.n1352 IREF.n1351 1.129
R7331 IREF.n1373 IREF.n1370 1.12765
R7332 IREF.n938 IREF.n937 1.11862
R7333 IREF.n1061 IREF.n1060 1.11862
R7334 IREF.n10 IREF.n9 0.9995
R7335 IREF.n18 IREF.n17 0.9995
R7336 IREF.n1296 IREF.n1295 0.915282
R7337 IREF.n1306 IREF.n1305 0.915282
R7338 IREF.n1317 IREF.n1316 0.915282
R7339 IREF.n1328 IREF.n1327 0.915282
R7340 IREF.n1339 IREF.n1338 0.915282
R7341 IREF.n1384 IREF.n37 0.886209
R7342 IREF.n430 IREF.n390 0.83975
R7343 IREF.n552 IREF.n131 0.83975
R7344 IREF.n1290 IREF.n40 0.83975
R7345 IREF.n1249 IREF.n1189 0.83975
R7346 IREF.n388 IREF.n160 0.81725
R7347 IREF.n257 IREF.n130 0.81725
R7348 IREF.n652 IREF.n651 0.81725
R7349 IREF.n783 IREF.n554 0.81725
R7350 IREF.n1117 IREF.n1116 0.809892
R7351 IREF.n1186 IREF.n785 0.809892
R7352 IREF.n1364 IREF.n1363 0.779178
R7353 IREF.n83 IREF.n82 0.75626
R7354 IREF.n1247 IREF.n1246 0.75626
R7355 IREF.n433 IREF.n432 0.75626
R7356 IREF.n502 IREF.n501 0.75626
R7357 IREF.n212 IREF.n211 0.756242
R7358 IREF.n324 IREF.n323 0.756242
R7359 IREF.n649 IREF.n648 0.756242
R7360 IREF.n724 IREF.n723 0.756242
R7361 IREF.n889 IREF.n816 0.752
R7362 IREF.n950 IREF.n949 0.752
R7363 IREF.n1115 IREF.n1114 0.752
R7364 IREF.n1071 IREF.n1053 0.752
R7365 IREF.n1014 IREF.n1013 0.71825
R7366 IREF.n971 IREF.n952 0.71825
R7367 IREF.n1118 IREF.n799 0.71825
R7368 IREF.n1185 IREF.n1184 0.71825
R7369 IREF.n96 IREF.n95 0.698
R7370 IREF.n1235 IREF.n1234 0.698
R7371 IREF.n385 IREF.n224 0.698
R7372 IREF.n312 IREF.n311 0.698
R7373 IREF.n447 IREF.n445 0.698
R7374 IREF.n515 IREF.n514 0.698
R7375 IREF.n656 IREF.n589 0.698
R7376 IREF.n780 IREF.n736 0.698
R7377 IREF.n1302 IREF.n1301 0.688348
R7378 IREF.n1312 IREF.n1311 0.688348
R7379 IREF.n1323 IREF.n1322 0.688348
R7380 IREF.n1334 IREF.n1333 0.688348
R7381 IREF.n1345 IREF.n1344 0.688348
R7382 IREF.n1164 IREF.n1163 0.673132
R7383 IREF.n1165 IREF.n1164 0.673132
R7384 IREF.n1122 IREF.n1121 0.673132
R7385 IREF.n1123 IREF.n1122 0.673132
R7386 IREF.n931 IREF.n930 0.673132
R7387 IREF.n932 IREF.n931 0.673132
R7388 IREF.n886 IREF.n885 0.673132
R7389 IREF.n887 IREF.n886 0.673132
R7390 IREF.n975 IREF.n974 0.673132
R7391 IREF.n974 IREF.n973 0.673132
R7392 IREF.n837 IREF.n836 0.673132
R7393 IREF.n838 IREF.n837 0.673132
R7394 IREF.n1075 IREF.n1074 0.673132
R7395 IREF.n1074 IREF.n1073 0.673132
R7396 IREF.n1038 IREF.n1037 0.673132
R7397 IREF.n1039 IREF.n1038 0.673132
R7398 IREF.n1297 IREF.n1296 0.655148
R7399 IREF.n1307 IREF.n1306 0.655148
R7400 IREF.n1318 IREF.n1317 0.655148
R7401 IREF.n1365 IREF.n1364 0.655148
R7402 IREF.n1329 IREF.n1328 0.655148
R7403 IREF.n1340 IREF.n1339 0.655148
R7404 IREF.n1295 IREF.n1294 0.63334
R7405 IREF.n1301 IREF.n1300 0.63334
R7406 IREF.n1300 IREF.n1299 0.63334
R7407 IREF.n1305 IREF.n1304 0.63334
R7408 IREF.n1311 IREF.n1310 0.63334
R7409 IREF.n1310 IREF.n1309 0.63334
R7410 IREF.n1316 IREF.n1315 0.63334
R7411 IREF.n1322 IREF.n1321 0.63334
R7412 IREF.n1321 IREF.n1320 0.63334
R7413 IREF.n1327 IREF.n1326 0.63334
R7414 IREF.n1333 IREF.n1332 0.63334
R7415 IREF.n1332 IREF.n1331 0.63334
R7416 IREF.n1338 IREF.n1337 0.63334
R7417 IREF.n1344 IREF.n1343 0.63334
R7418 IREF.n1343 IREF.n1342 0.63334
R7419 IREF.n1294 IREF.n1293 0.63225
R7420 IREF.n1298 IREF.n1297 0.63225
R7421 IREF.n1304 IREF.n1303 0.63225
R7422 IREF.n1308 IREF.n1307 0.63225
R7423 IREF.n1315 IREF.n1314 0.63225
R7424 IREF.n1319 IREF.n1318 0.63225
R7425 IREF.n1366 IREF.n1365 0.63225
R7426 IREF.n1326 IREF.n1325 0.63225
R7427 IREF.n1330 IREF.n1329 0.63225
R7428 IREF.n1337 IREF.n1336 0.63225
R7429 IREF.n1341 IREF.n1340 0.63225
R7430 IREF.n1381 IREF.n1380 0.622055
R7431 IREF.n1292 IREF.n38 0.602344
R7432 IREF.n1291 IREF.n39 0.571818
R7433 IREF.n1188 IREF.n784 0.571818
R7434 IREF.n1335 IREF.n1324 0.467527
R7435 IREF.n1170 IREF.n1169 0.45279
R7436 IREF.n959 IREF.n958 0.45279
R7437 IREF.n870 IREF.n869 0.430924
R7438 IREF.n1022 IREF.n1021 0.430924
R7439 IREF.n940 IREF.n939 0.394842
R7440 IREF.n920 IREF.n856 0.394842
R7441 IREF.n899 IREF.n898 0.394842
R7442 IREF.n875 IREF.n873 0.394842
R7443 IREF.n1063 IREF.n1062 0.394842
R7444 IREF.n1086 IREF.n1085 0.394842
R7445 IREF.n1105 IREF.n1104 0.394842
R7446 IREF.n1027 IREF.n1020 0.394842
R7447 IREF.n945 IREF.n933 0.381816
R7448 IREF.n914 IREF.n913 0.381816
R7449 IREF.n894 IREF.n892 0.381816
R7450 IREF.n1068 IREF.n1067 0.381816
R7451 IREF.n1091 IREF.n1047 0.381816
R7452 IREF.n1110 IREF.n1040 0.381816
R7453 IREF.n1180 IREF.n1166 0.379447
R7454 IREF.n1174 IREF.n1173 0.379447
R7455 IREF.n1147 IREF.n1146 0.379447
R7456 IREF.n1153 IREF.n790 0.379447
R7457 IREF.n1156 IREF.n788 0.379447
R7458 IREF.n1129 IREF.n1128 0.379447
R7459 IREF.n1134 IREF.n1133 0.379447
R7460 IREF.n1140 IREF.n794 0.379447
R7461 IREF.n808 IREF.n807 0.379447
R7462 IREF.n813 IREF.n812 0.379447
R7463 IREF.n968 IREF.n967 0.379447
R7464 IREF.n963 IREF.n962 0.379447
R7465 IREF.n991 IREF.n990 0.379447
R7466 IREF.n986 IREF.n985 0.379447
R7467 IREF.n981 IREF.n980 0.379447
R7468 IREF.n1009 IREF.n839 0.379447
R7469 IREF.n1003 IREF.n1002 0.379447
R7470 IREF.n998 IREF.n997 0.379447
R7471 IREF.n826 IREF.n821 0.379447
R7472 IREF.n829 IREF.n819 0.379447
R7473 IREF.n1378 IREF.n1377 0.379447
R7474 IREF.n1372 IREF.n1369 0.379447
R7475 IREF.n1360 IREF.n1348 0.379447
R7476 IREF.n1354 IREF.n1353 0.378263
R7477 IREF.n71 IREF.n50 0.375125
R7478 IREF.n105 IREF.n104 0.375125
R7479 IREF.n125 IREF.n121 0.375125
R7480 IREF.n1206 IREF.n1205 0.375125
R7481 IREF.n192 IREF.n171 0.375125
R7482 IREF.n369 IREF.n230 0.375125
R7483 IREF.n342 IREF.n251 0.375125
R7484 IREF.n296 IREF.n295 0.375125
R7485 IREF.n417 IREF.n399 0.375125
R7486 IREF.n462 IREF.n153 0.375125
R7487 IREF.n490 IREF.n141 0.375125
R7488 IREF.n524 IREF.n523 0.375125
R7489 IREF.n420 IREF.n401 0.375125
R7490 IREF.n460 IREF.n459 0.375125
R7491 IREF.n488 IREF.n487 0.375125
R7492 IREF.n540 IREF.n519 0.375125
R7493 IREF.n622 IREF.n596 0.375125
R7494 IREF.n675 IREF.n581 0.375125
R7495 IREF.n704 IREF.n565 0.375125
R7496 IREF.n764 IREF.n742 0.375125
R7497 IREF.n69 IREF.n68 0.375125
R7498 IREF.n1278 IREF.n100 0.375125
R7499 IREF.n1257 IREF.n1256 0.375125
R7500 IREF.n1222 IREF.n1203 0.375125
R7501 IREF.n876 IREF.n868 0.375125
R7502 IREF.n897 IREF.n861 0.375125
R7503 IREF.n919 IREF.n918 0.375125
R7504 IREF.n938 IREF.n934 0.375125
R7505 IREF.n1026 IREF.n1025 0.375125
R7506 IREF.n1103 IREF.n1041 0.375125
R7507 IREF.n1084 IREF.n1048 0.375125
R7508 IREF.n1061 IREF.n1058 0.375125
R7509 IREF.n64 IREF.n55 0.36275
R7510 IREF.n102 IREF.n98 0.36275
R7511 IREF.n119 IREF.n118 0.36275
R7512 IREF.n1201 IREF.n1200 0.36275
R7513 IREF.n183 IREF.n175 0.36275
R7514 IREF.n377 IREF.n225 0.36275
R7515 IREF.n351 IREF.n246 0.36275
R7516 IREF.n304 IREF.n303 0.36275
R7517 IREF.n415 IREF.n403 0.36275
R7518 IREF.n455 IREF.n158 0.36275
R7519 IREF.n483 IREF.n146 0.36275
R7520 IREF.n521 IREF.n517 0.36275
R7521 IREF.n413 IREF.n411 0.36275
R7522 IREF.n452 IREF.n156 0.36275
R7523 IREF.n480 IREF.n144 0.36275
R7524 IREF.n546 IREF.n545 0.36275
R7525 IREF.n612 IREF.n600 0.36275
R7526 IREF.n665 IREF.n585 0.36275
R7527 IREF.n695 IREF.n569 0.36275
R7528 IREF.n772 IREF.n737 0.36275
R7529 IREF.n61 IREF.n53 0.36275
R7530 IREF.n1284 IREF.n1283 0.36275
R7531 IREF.n1263 IREF.n1262 0.36275
R7532 IREF.n1227 IREF.n1199 0.36275
R7533 IREF.n895 IREF.n863 0.36275
R7534 IREF.n912 IREF.n857 0.36275
R7535 IREF.n944 IREF.n943 0.36275
R7536 IREF.n1109 IREF.n1108 0.36275
R7537 IREF.n1090 IREF.n1089 0.36275
R7538 IREF.n1066 IREF.n1056 0.36275
R7539 IREF.n84 IREF.n44 0.3605
R7540 IREF.n91 IREF.n90 0.3605
R7541 IREF.n1242 IREF.n1192 0.3605
R7542 IREF.n1240 IREF.n1194 0.3605
R7543 IREF.n213 IREF.n165 0.3605
R7544 IREF.n220 IREF.n219 0.3605
R7545 IREF.n319 IREF.n259 0.3605
R7546 IREF.n317 IREF.n261 0.3605
R7547 IREF.n186 IREF.n177 0.3605
R7548 IREF.n195 IREF.n173 0.3605
R7549 IREF.n206 IREF.n169 0.3605
R7550 IREF.n381 IREF.n380 0.3605
R7551 IREF.n373 IREF.n372 0.3605
R7552 IREF.n365 IREF.n364 0.3605
R7553 IREF.n348 IREF.n248 0.3605
R7554 IREF.n339 IREF.n249 0.3605
R7555 IREF.n329 IREF.n253 0.3605
R7556 IREF.n307 IREF.n267 0.3605
R7557 IREF.n299 IREF.n272 0.3605
R7558 IREF.n291 IREF.n277 0.3605
R7559 IREF.n434 IREF.n393 0.3605
R7560 IREF.n441 IREF.n440 0.3605
R7561 IREF.n503 IREF.n135 0.3605
R7562 IREF.n510 IREF.n509 0.3605
R7563 IREF.n644 IREF.n633 0.3605
R7564 IREF.n642 IREF.n635 0.3605
R7565 IREF.n725 IREF.n559 0.3605
R7566 IREF.n732 IREF.n731 0.3605
R7567 IREF.n608 IREF.n607 0.3605
R7568 IREF.n617 IREF.n616 0.3605
R7569 IREF.n628 IREF.n627 0.3605
R7570 IREF.n661 IREF.n660 0.3605
R7571 IREF.n670 IREF.n669 0.3605
R7572 IREF.n681 IREF.n680 0.3605
R7573 IREF.n698 IREF.n571 0.3605
R7574 IREF.n707 IREF.n567 0.3605
R7575 IREF.n718 IREF.n563 0.3605
R7576 IREF.n776 IREF.n775 0.3605
R7577 IREF.n768 IREF.n767 0.3605
R7578 IREF.n760 IREF.n759 0.3605
R7579 IREF.n825 IREF.n824 0.3605
R7580 IREF.n831 IREF.n830 0.3605
R7581 IREF.n1008 IREF.n1007 0.3605
R7582 IREF.n1001 IREF.n840 0.3605
R7583 IREF.n999 IREF.n842 0.3605
R7584 IREF.n989 IREF.n845 0.3605
R7585 IREF.n987 IREF.n847 0.3605
R7586 IREF.n982 IREF.n850 0.3605
R7587 IREF.n969 IREF.n954 0.3605
R7588 IREF.n964 IREF.n957 0.3605
R7589 IREF.n806 IREF.n803 0.3605
R7590 IREF.n811 IREF.n801 0.3605
R7591 IREF.n1127 IREF.n797 0.3605
R7592 IREF.n1132 IREF.n795 0.3605
R7593 IREF.n1139 IREF.n1138 0.3605
R7594 IREF.n1145 IREF.n791 0.3605
R7595 IREF.n1152 IREF.n1151 0.3605
R7596 IREF.n1158 IREF.n1157 0.3605
R7597 IREF.n1179 IREF.n1178 0.3605
R7598 IREF.n1172 IREF.n1167 0.3605
R7599 IREF.n1359 IREF.n1358 0.3605
R7600 IREF.n1379 IREF.n1368 0.3605
R7601 IREF.n1374 IREF.n1373 0.3605
R7602 IREF.n1352 IREF.n1349 0.359375
R7603 IREF.n937 IREF.n936 0.348488
R7604 IREF.n1060 IREF.n1059 0.348488
R7605 IREF.n805 IREF.n804 0.327481
R7606 IREF.n823 IREF.n822 0.327481
R7607 IREF.n1351 IREF.n1350 0.32675
R7608 IREF.n1371 IREF.n1370 0.324133
R7609 IREF.n1346 IREF.n1335 0.307291
R7610 IREF.n923 IREF.n854 0.302474
R7611 IREF.n905 IREF.n860 0.302474
R7612 IREF.n880 IREF.n879 0.302474
R7613 IREF.n1081 IREF.n1080 0.302474
R7614 IREF.n1100 IREF.n1099 0.302474
R7615 IREF.n1030 IREF.n1018 0.302474
R7616 IREF.n1324 IREF.n1313 0.301209
R7617 IREF.n74 IREF.n73 0.287375
R7618 IREF.n110 IREF.n109 0.287375
R7619 IREF.n128 IREF.n127 0.287375
R7620 IREF.n1211 IREF.n1210 0.287375
R7621 IREF.n203 IREF.n202 0.287375
R7622 IREF.n241 IREF.n235 0.287375
R7623 IREF.n333 IREF.n255 0.287375
R7624 IREF.n288 IREF.n287 0.287375
R7625 IREF.n426 IREF.n425 0.287375
R7626 IREF.n465 IREF.n464 0.287375
R7627 IREF.n493 IREF.n492 0.287375
R7628 IREF.n529 IREF.n528 0.287375
R7629 IREF.n421 IREF.n397 0.287375
R7630 IREF.n468 IREF.n467 0.287375
R7631 IREF.n496 IREF.n495 0.287375
R7632 IREF.n535 IREF.n526 0.287375
R7633 IREF.n624 IREF.n592 0.287375
R7634 IREF.n677 IREF.n577 0.287375
R7635 IREF.n715 IREF.n714 0.287375
R7636 IREF.n753 IREF.n747 0.287375
R7637 IREF.n77 IREF.n76 0.287375
R7638 IREF.n1273 IREF.n107 0.287375
R7639 IREF.n1251 IREF.n123 0.287375
R7640 IREF.n1217 IREF.n1208 0.287375
R7641 IREF.n878 IREF.n866 0.287375
R7642 IREF.n904 IREF.n903 0.287375
R7643 IREF.n925 IREF.n924 0.287375
R7644 IREF.n1032 IREF.n1031 0.287375
R7645 IREF.n1098 IREF.n1044 0.287375
R7646 IREF.n1079 IREF.n1051 0.287375
R7647 IREF.n1302 IREF.n1298 0.254694
R7648 IREF.n1312 IREF.n1308 0.254694
R7649 IREF.n1323 IREF.n1319 0.254694
R7650 IREF.n1381 IREF.n1366 0.254694
R7651 IREF.n1334 IREF.n1330 0.254694
R7652 IREF.n1345 IREF.n1341 0.254694
R7653 IREF.n213 IREF.n212 0.208888
R7654 IREF.n323 IREF.n259 0.208888
R7655 IREF.n648 IREF.n633 0.208888
R7656 IREF.n725 IREF.n724 0.208888
R7657 IREF.n84 IREF.n83 0.20887
R7658 IREF.n1246 IREF.n1192 0.20887
R7659 IREF.n434 IREF.n433 0.20887
R7660 IREF.n503 IREF.n502 0.20887
R7661 IREF.n993 IREF.n845 0.208099
R7662 IREF.n1145 IREF.n1144 0.208099
R7663 IREF.n1380 IREF.n1379 0.208099
R7664 IREF.n1183 IREF.n1182 0.147342
R7665 IREF.n1176 IREF.n1166 0.147342
R7666 IREF.n1173 IREF.n1168 0.147342
R7667 IREF.n1149 IREF.n1147 0.147342
R7668 IREF.n1154 IREF.n1153 0.147342
R7669 IREF.n1160 IREF.n788 0.147342
R7670 IREF.n1125 IREF.n1124 0.147342
R7671 IREF.n1130 IREF.n1129 0.147342
R7672 IREF.n1136 IREF.n1134 0.147342
R7673 IREF.n1141 IREF.n1140 0.147342
R7674 IREF.n809 IREF.n808 0.147342
R7675 IREF.n814 IREF.n813 0.147342
R7676 IREF.n946 IREF.n945 0.147342
R7677 IREF.n941 IREF.n940 0.147342
R7678 IREF.n913 IREF.n858 0.147342
R7679 IREF.n916 IREF.n856 0.147342
R7680 IREF.n923 IREF.n922 0.147342
R7681 IREF.n927 IREF.n854 0.147342
R7682 IREF.n892 IREF.n891 0.147342
R7683 IREF.n898 IREF.n862 0.147342
R7684 IREF.n901 IREF.n860 0.147342
R7685 IREF.n906 IREF.n905 0.147342
R7686 IREF.n873 IREF.n872 0.147342
R7687 IREF.n879 IREF.n867 0.147342
R7688 IREF.n881 IREF.n880 0.147342
R7689 IREF.n972 IREF.n953 0.147342
R7690 IREF.n967 IREF.n966 0.147342
R7691 IREF.n962 IREF.n961 0.147342
R7692 IREF.n990 IREF.n846 0.147342
R7693 IREF.n985 IREF.n984 0.147342
R7694 IREF.n980 IREF.n979 0.147342
R7695 IREF.n1012 IREF.n1011 0.147342
R7696 IREF.n1005 IREF.n839 0.147342
R7697 IREF.n1002 IREF.n841 0.147342
R7698 IREF.n997 IREF.n996 0.147342
R7699 IREF.n827 IREF.n826 0.147342
R7700 IREF.n833 IREF.n819 0.147342
R7701 IREF.n1069 IREF.n1068 0.147342
R7702 IREF.n1064 IREF.n1063 0.147342
R7703 IREF.n1092 IREF.n1091 0.147342
R7704 IREF.n1087 IREF.n1086 0.147342
R7705 IREF.n1082 IREF.n1081 0.147342
R7706 IREF.n1080 IREF.n1052 0.147342
R7707 IREF.n1111 IREF.n1110 0.147342
R7708 IREF.n1106 IREF.n1105 0.147342
R7709 IREF.n1101 IREF.n1100 0.147342
R7710 IREF.n1099 IREF.n1045 0.147342
R7711 IREF.n1023 IREF.n1020 0.147342
R7712 IREF.n1030 IREF.n1029 0.147342
R7713 IREF.n1034 IREF.n1018 0.147342
R7714 IREF.n1378 IREF.n1367 0.147342
R7715 IREF.n1377 IREF.n1376 0.147342
R7716 IREF.n1376 IREF.n1369 0.147342
R7717 IREF.n1372 IREF.n1371 0.147342
R7718 IREF.n1356 IREF.n1354 0.147342
R7719 IREF.n1361 IREF.n1360 0.147342
R7720 IREF.n1353 IREF.n1350 0.143789
R7721 IREF.n1181 IREF.n1180 0.142605
R7722 IREF.n1175 IREF.n1174 0.142605
R7723 IREF.n1146 IREF.n792 0.142605
R7724 IREF.n1148 IREF.n790 0.142605
R7725 IREF.n1156 IREF.n1155 0.142605
R7726 IREF.n1162 IREF.n1161 0.142605
R7727 IREF.n1128 IREF.n798 0.142605
R7728 IREF.n1133 IREF.n796 0.142605
R7729 IREF.n1135 IREF.n794 0.142605
R7730 IREF.n807 IREF.n804 0.142605
R7731 IREF.n812 IREF.n802 0.142605
R7732 IREF.n1120 IREF.n800 0.142605
R7733 IREF.n968 IREF.n955 0.142605
R7734 IREF.n963 IREF.n956 0.142605
R7735 IREF.n992 IREF.n991 0.142605
R7736 IREF.n986 IREF.n848 0.142605
R7737 IREF.n981 IREF.n849 0.142605
R7738 IREF.n976 IREF.n851 0.142605
R7739 IREF.n1010 IREF.n1009 0.142605
R7740 IREF.n1004 IREF.n1003 0.142605
R7741 IREF.n998 IREF.n843 0.142605
R7742 IREF.n822 IREF.n821 0.142605
R7743 IREF.n829 IREF.n828 0.142605
R7744 IREF.n835 IREF.n834 0.142605
R7745 IREF.n1355 IREF.n1348 0.142605
R7746 IREF.n33 IREF.n29 0.14
R7747 IREF.n36 IREF.n29 0.14
R7748 IREF.n57 IREF.n55 0.14
R7749 IREF.n65 IREF.n64 0.14
R7750 IREF.n65 IREF.n50 0.14
R7751 IREF.n72 IREF.n71 0.14
R7752 IREF.n74 IREF.n72 0.14
R7753 IREF.n73 IREF.n46 0.14
R7754 IREF.n82 IREF.n46 0.14
R7755 IREF.n89 IREF.n44 0.14
R7756 IREF.n90 IREF.n89 0.14
R7757 IREF.n91 IREF.n42 0.14
R7758 IREF.n95 IREF.n42 0.14
R7759 IREF.n97 IREF.n96 0.14
R7760 IREF.n98 IREF.n97 0.14
R7761 IREF.n103 IREF.n102 0.14
R7762 IREF.n104 IREF.n103 0.14
R7763 IREF.n108 IREF.n105 0.14
R7764 IREF.n109 IREF.n108 0.14
R7765 IREF.n114 IREF.n110 0.14
R7766 IREF.n1269 IREF.n114 0.14
R7767 IREF.n1268 IREF.n115 0.14
R7768 IREF.n118 IREF.n115 0.14
R7769 IREF.n120 IREF.n119 0.14
R7770 IREF.n121 IREF.n120 0.14
R7771 IREF.n126 IREF.n125 0.14
R7772 IREF.n127 IREF.n126 0.14
R7773 IREF.n1191 IREF.n128 0.14
R7774 IREF.n1247 IREF.n1191 0.14
R7775 IREF.n1242 IREF.n1241 0.14
R7776 IREF.n1241 IREF.n1240 0.14
R7777 IREF.n1236 IREF.n1194 0.14
R7778 IREF.n1236 IREF.n1235 0.14
R7779 IREF.n1234 IREF.n1197 0.14
R7780 IREF.n1200 IREF.n1197 0.14
R7781 IREF.n1204 IREF.n1201 0.14
R7782 IREF.n1205 IREF.n1204 0.14
R7783 IREF.n1209 IREF.n1206 0.14
R7784 IREF.n1210 IREF.n1209 0.14
R7785 IREF.n1214 IREF.n1211 0.14
R7786 IREF.n183 IREF.n182 0.14
R7787 IREF.n191 IREF.n175 0.14
R7788 IREF.n192 IREF.n191 0.14
R7789 IREF.n201 IREF.n171 0.14
R7790 IREF.n202 IREF.n201 0.14
R7791 IREF.n203 IREF.n167 0.14
R7792 IREF.n211 IREF.n167 0.14
R7793 IREF.n218 IREF.n165 0.14
R7794 IREF.n219 IREF.n218 0.14
R7795 IREF.n220 IREF.n163 0.14
R7796 IREF.n224 IREF.n163 0.14
R7797 IREF.n385 IREF.n384 0.14
R7798 IREF.n384 IREF.n225 0.14
R7799 IREF.n377 IREF.n376 0.14
R7800 IREF.n376 IREF.n230 0.14
R7801 IREF.n369 IREF.n368 0.14
R7802 IREF.n368 IREF.n235 0.14
R7803 IREF.n361 IREF.n241 0.14
R7804 IREF.n361 IREF.n360 0.14
R7805 IREF.n352 IREF.n242 0.14
R7806 IREF.n352 IREF.n351 0.14
R7807 IREF.n343 IREF.n246 0.14
R7808 IREF.n343 IREF.n342 0.14
R7809 IREF.n334 IREF.n251 0.14
R7810 IREF.n334 IREF.n333 0.14
R7811 IREF.n258 IREF.n255 0.14
R7812 IREF.n324 IREF.n258 0.14
R7813 IREF.n319 IREF.n318 0.14
R7814 IREF.n318 IREF.n317 0.14
R7815 IREF.n313 IREF.n261 0.14
R7816 IREF.n313 IREF.n312 0.14
R7817 IREF.n311 IREF.n264 0.14
R7818 IREF.n304 IREF.n264 0.14
R7819 IREF.n303 IREF.n270 0.14
R7820 IREF.n296 IREF.n270 0.14
R7821 IREF.n295 IREF.n275 0.14
R7822 IREF.n288 IREF.n275 0.14
R7823 IREF.n287 IREF.n286 0.14
R7824 IREF.n187 IREF.n186 0.14
R7825 IREF.n187 IREF.n173 0.14
R7826 IREF.n196 IREF.n195 0.14
R7827 IREF.n196 IREF.n169 0.14
R7828 IREF.n207 IREF.n206 0.14
R7829 IREF.n207 IREF.n160 0.14
R7830 IREF.n387 IREF.n161 0.14
R7831 IREF.n381 IREF.n161 0.14
R7832 IREF.n380 IREF.n228 0.14
R7833 IREF.n373 IREF.n228 0.14
R7834 IREF.n372 IREF.n233 0.14
R7835 IREF.n365 IREF.n233 0.14
R7836 IREF.n364 IREF.n238 0.14
R7837 IREF.n358 IREF.n238 0.14
R7838 IREF.n357 IREF.n244 0.14
R7839 IREF.n248 IREF.n244 0.14
R7840 IREF.n348 IREF.n347 0.14
R7841 IREF.n347 IREF.n249 0.14
R7842 IREF.n339 IREF.n338 0.14
R7843 IREF.n338 IREF.n253 0.14
R7844 IREF.n329 IREF.n328 0.14
R7845 IREF.n328 IREF.n257 0.14
R7846 IREF.n308 IREF.n265 0.14
R7847 IREF.n308 IREF.n307 0.14
R7848 IREF.n300 IREF.n267 0.14
R7849 IREF.n300 IREF.n299 0.14
R7850 IREF.n292 IREF.n272 0.14
R7851 IREF.n292 IREF.n291 0.14
R7852 IREF.n283 IREF.n277 0.14
R7853 IREF.n408 IREF.n403 0.14
R7854 IREF.n416 IREF.n415 0.14
R7855 IREF.n417 IREF.n416 0.14
R7856 IREF.n424 IREF.n399 0.14
R7857 IREF.n425 IREF.n424 0.14
R7858 IREF.n426 IREF.n395 0.14
R7859 IREF.n432 IREF.n395 0.14
R7860 IREF.n439 IREF.n393 0.14
R7861 IREF.n440 IREF.n439 0.14
R7862 IREF.n441 IREF.n391 0.14
R7863 IREF.n445 IREF.n391 0.14
R7864 IREF.n447 IREF.n446 0.14
R7865 IREF.n446 IREF.n158 0.14
R7866 IREF.n456 IREF.n455 0.14
R7867 IREF.n456 IREF.n153 0.14
R7868 IREF.n463 IREF.n462 0.14
R7869 IREF.n465 IREF.n463 0.14
R7870 IREF.n464 IREF.n149 0.14
R7871 IREF.n473 IREF.n149 0.14
R7872 IREF.n475 IREF.n474 0.14
R7873 IREF.n474 IREF.n146 0.14
R7874 IREF.n484 IREF.n483 0.14
R7875 IREF.n484 IREF.n141 0.14
R7876 IREF.n491 IREF.n490 0.14
R7877 IREF.n493 IREF.n491 0.14
R7878 IREF.n492 IREF.n137 0.14
R7879 IREF.n501 IREF.n137 0.14
R7880 IREF.n508 IREF.n135 0.14
R7881 IREF.n509 IREF.n508 0.14
R7882 IREF.n510 IREF.n133 0.14
R7883 IREF.n514 IREF.n133 0.14
R7884 IREF.n516 IREF.n515 0.14
R7885 IREF.n517 IREF.n516 0.14
R7886 IREF.n522 IREF.n521 0.14
R7887 IREF.n523 IREF.n522 0.14
R7888 IREF.n527 IREF.n524 0.14
R7889 IREF.n528 IREF.n527 0.14
R7890 IREF.n532 IREF.n529 0.14
R7891 IREF.n411 IREF.n410 0.14
R7892 IREF.n413 IREF.n412 0.14
R7893 IREF.n412 IREF.n401 0.14
R7894 IREF.n422 IREF.n420 0.14
R7895 IREF.n422 IREF.n421 0.14
R7896 IREF.n429 IREF.n397 0.14
R7897 IREF.n430 IREF.n429 0.14
R7898 IREF.n451 IREF.n450 0.14
R7899 IREF.n452 IREF.n451 0.14
R7900 IREF.n458 IREF.n156 0.14
R7901 IREF.n459 IREF.n458 0.14
R7902 IREF.n460 IREF.n151 0.14
R7903 IREF.n467 IREF.n151 0.14
R7904 IREF.n469 IREF.n468 0.14
R7905 IREF.n469 IREF.n148 0.14
R7906 IREF.n479 IREF.n478 0.14
R7907 IREF.n480 IREF.n479 0.14
R7908 IREF.n486 IREF.n144 0.14
R7909 IREF.n487 IREF.n486 0.14
R7910 IREF.n488 IREF.n139 0.14
R7911 IREF.n495 IREF.n139 0.14
R7912 IREF.n497 IREF.n496 0.14
R7913 IREF.n497 IREF.n131 0.14
R7914 IREF.n551 IREF.n132 0.14
R7915 IREF.n546 IREF.n132 0.14
R7916 IREF.n545 IREF.n544 0.14
R7917 IREF.n544 IREF.n519 0.14
R7918 IREF.n540 IREF.n539 0.14
R7919 IREF.n539 IREF.n526 0.14
R7920 IREF.n535 IREF.n534 0.14
R7921 IREF.n604 IREF.n600 0.14
R7922 IREF.n613 IREF.n612 0.14
R7923 IREF.n613 IREF.n596 0.14
R7924 IREF.n623 IREF.n622 0.14
R7925 IREF.n624 IREF.n623 0.14
R7926 IREF.n632 IREF.n592 0.14
R7927 IREF.n649 IREF.n632 0.14
R7928 IREF.n644 IREF.n643 0.14
R7929 IREF.n643 IREF.n642 0.14
R7930 IREF.n638 IREF.n635 0.14
R7931 IREF.n638 IREF.n589 0.14
R7932 IREF.n657 IREF.n656 0.14
R7933 IREF.n657 IREF.n585 0.14
R7934 IREF.n666 IREF.n665 0.14
R7935 IREF.n666 IREF.n581 0.14
R7936 IREF.n676 IREF.n675 0.14
R7937 IREF.n677 IREF.n676 0.14
R7938 IREF.n685 IREF.n577 0.14
R7939 IREF.n686 IREF.n685 0.14
R7940 IREF.n694 IREF.n573 0.14
R7941 IREF.n695 IREF.n694 0.14
R7942 IREF.n703 IREF.n569 0.14
R7943 IREF.n704 IREF.n703 0.14
R7944 IREF.n713 IREF.n565 0.14
R7945 IREF.n714 IREF.n713 0.14
R7946 IREF.n715 IREF.n561 0.14
R7947 IREF.n723 IREF.n561 0.14
R7948 IREF.n730 IREF.n559 0.14
R7949 IREF.n731 IREF.n730 0.14
R7950 IREF.n732 IREF.n557 0.14
R7951 IREF.n736 IREF.n557 0.14
R7952 IREF.n780 IREF.n779 0.14
R7953 IREF.n779 IREF.n737 0.14
R7954 IREF.n772 IREF.n771 0.14
R7955 IREF.n771 IREF.n742 0.14
R7956 IREF.n764 IREF.n763 0.14
R7957 IREF.n763 IREF.n747 0.14
R7958 IREF.n756 IREF.n753 0.14
R7959 IREF.n608 IREF.n598 0.14
R7960 IREF.n616 IREF.n598 0.14
R7961 IREF.n617 IREF.n594 0.14
R7962 IREF.n627 IREF.n594 0.14
R7963 IREF.n628 IREF.n590 0.14
R7964 IREF.n651 IREF.n590 0.14
R7965 IREF.n653 IREF.n587 0.14
R7966 IREF.n660 IREF.n587 0.14
R7967 IREF.n661 IREF.n583 0.14
R7968 IREF.n669 IREF.n583 0.14
R7969 IREF.n670 IREF.n579 0.14
R7970 IREF.n680 IREF.n579 0.14
R7971 IREF.n681 IREF.n575 0.14
R7972 IREF.n688 IREF.n575 0.14
R7973 IREF.n690 IREF.n689 0.14
R7974 IREF.n690 IREF.n571 0.14
R7975 IREF.n699 IREF.n698 0.14
R7976 IREF.n699 IREF.n567 0.14
R7977 IREF.n708 IREF.n707 0.14
R7978 IREF.n708 IREF.n563 0.14
R7979 IREF.n719 IREF.n718 0.14
R7980 IREF.n719 IREF.n554 0.14
R7981 IREF.n782 IREF.n555 0.14
R7982 IREF.n776 IREF.n555 0.14
R7983 IREF.n775 IREF.n740 0.14
R7984 IREF.n768 IREF.n740 0.14
R7985 IREF.n767 IREF.n745 0.14
R7986 IREF.n760 IREF.n745 0.14
R7987 IREF.n759 IREF.n750 0.14
R7988 IREF.n61 IREF.n60 0.14
R7989 IREF.n67 IREF.n53 0.14
R7990 IREF.n68 IREF.n67 0.14
R7991 IREF.n69 IREF.n48 0.14
R7992 IREF.n76 IREF.n48 0.14
R7993 IREF.n78 IREF.n77 0.14
R7994 IREF.n78 IREF.n40 0.14
R7995 IREF.n1289 IREF.n41 0.14
R7996 IREF.n1284 IREF.n41 0.14
R7997 IREF.n1283 IREF.n1282 0.14
R7998 IREF.n1282 IREF.n100 0.14
R7999 IREF.n1278 IREF.n1277 0.14
R8000 IREF.n1277 IREF.n107 0.14
R8001 IREF.n1273 IREF.n1272 0.14
R8002 IREF.n1272 IREF.n1271 0.14
R8003 IREF.n1264 IREF.n112 0.14
R8004 IREF.n1264 IREF.n1263 0.14
R8005 IREF.n1262 IREF.n117 0.14
R8006 IREF.n1257 IREF.n117 0.14
R8007 IREF.n1256 IREF.n1255 0.14
R8008 IREF.n1255 IREF.n123 0.14
R8009 IREF.n1251 IREF.n1250 0.14
R8010 IREF.n1250 IREF.n1249 0.14
R8011 IREF.n1232 IREF.n1231 0.14
R8012 IREF.n1231 IREF.n1199 0.14
R8013 IREF.n1227 IREF.n1226 0.14
R8014 IREF.n1226 IREF.n1203 0.14
R8015 IREF.n1222 IREF.n1221 0.14
R8016 IREF.n1221 IREF.n1208 0.14
R8017 IREF.n1217 IREF.n1216 0.14
R8018 IREF.n871 IREF.n868 0.14
R8019 IREF.n877 IREF.n876 0.14
R8020 IREF.n878 IREF.n877 0.14
R8021 IREF.n882 IREF.n866 0.14
R8022 IREF.n883 IREF.n882 0.14
R8023 IREF.n890 IREF.n889 0.14
R8024 IREF.n890 IREF.n863 0.14
R8025 IREF.n896 IREF.n895 0.14
R8026 IREF.n897 IREF.n896 0.14
R8027 IREF.n902 IREF.n861 0.14
R8028 IREF.n903 IREF.n902 0.14
R8029 IREF.n904 IREF.n859 0.14
R8030 IREF.n908 IREF.n859 0.14
R8031 IREF.n911 IREF.n910 0.14
R8032 IREF.n912 IREF.n911 0.14
R8033 IREF.n917 IREF.n857 0.14
R8034 IREF.n918 IREF.n917 0.14
R8035 IREF.n919 IREF.n855 0.14
R8036 IREF.n924 IREF.n855 0.14
R8037 IREF.n926 IREF.n925 0.14
R8038 IREF.n926 IREF.n852 0.14
R8039 IREF.n949 IREF.n853 0.14
R8040 IREF.n944 IREF.n853 0.14
R8041 IREF.n943 IREF.n942 0.14
R8042 IREF.n942 IREF.n934 0.14
R8043 IREF.n825 IREF.n820 0.14
R8044 IREF.n830 IREF.n820 0.14
R8045 IREF.n832 IREF.n831 0.14
R8046 IREF.n832 IREF.n817 0.14
R8047 IREF.n1013 IREF.n818 0.14
R8048 IREF.n1008 IREF.n818 0.14
R8049 IREF.n1007 IREF.n1006 0.14
R8050 IREF.n1006 IREF.n840 0.14
R8051 IREF.n1001 IREF.n1000 0.14
R8052 IREF.n1000 IREF.n999 0.14
R8053 IREF.n995 IREF.n842 0.14
R8054 IREF.n995 IREF.n994 0.14
R8055 IREF.n989 IREF.n988 0.14
R8056 IREF.n988 IREF.n987 0.14
R8057 IREF.n983 IREF.n847 0.14
R8058 IREF.n983 IREF.n982 0.14
R8059 IREF.n978 IREF.n850 0.14
R8060 IREF.n978 IREF.n977 0.14
R8061 IREF.n971 IREF.n970 0.14
R8062 IREF.n970 IREF.n969 0.14
R8063 IREF.n965 IREF.n954 0.14
R8064 IREF.n965 IREF.n964 0.14
R8065 IREF.n960 IREF.n957 0.14
R8066 IREF.n1025 IREF.n1024 0.14
R8067 IREF.n1026 IREF.n1019 0.14
R8068 IREF.n1031 IREF.n1019 0.14
R8069 IREF.n1033 IREF.n1032 0.14
R8070 IREF.n1033 IREF.n1016 0.14
R8071 IREF.n1114 IREF.n1017 0.14
R8072 IREF.n1109 IREF.n1017 0.14
R8073 IREF.n1108 IREF.n1107 0.14
R8074 IREF.n1107 IREF.n1041 0.14
R8075 IREF.n1103 IREF.n1102 0.14
R8076 IREF.n1102 IREF.n1044 0.14
R8077 IREF.n1098 IREF.n1097 0.14
R8078 IREF.n1097 IREF.n1096 0.14
R8079 IREF.n1094 IREF.n1046 0.14
R8080 IREF.n1090 IREF.n1046 0.14
R8081 IREF.n1089 IREF.n1088 0.14
R8082 IREF.n1088 IREF.n1048 0.14
R8083 IREF.n1084 IREF.n1083 0.14
R8084 IREF.n1083 IREF.n1051 0.14
R8085 IREF.n1079 IREF.n1078 0.14
R8086 IREF.n1078 IREF.n1077 0.14
R8087 IREF.n1071 IREF.n1070 0.14
R8088 IREF.n1070 IREF.n1056 0.14
R8089 IREF.n1066 IREF.n1065 0.14
R8090 IREF.n1065 IREF.n1058 0.14
R8091 IREF.n810 IREF.n803 0.14
R8092 IREF.n811 IREF.n810 0.14
R8093 IREF.n815 IREF.n801 0.14
R8094 IREF.n1119 IREF.n815 0.14
R8095 IREF.n1126 IREF.n799 0.14
R8096 IREF.n1127 IREF.n1126 0.14
R8097 IREF.n1131 IREF.n797 0.14
R8098 IREF.n1132 IREF.n1131 0.14
R8099 IREF.n1137 IREF.n795 0.14
R8100 IREF.n1138 IREF.n1137 0.14
R8101 IREF.n1139 IREF.n793 0.14
R8102 IREF.n1143 IREF.n793 0.14
R8103 IREF.n1150 IREF.n791 0.14
R8104 IREF.n1151 IREF.n1150 0.14
R8105 IREF.n1152 IREF.n789 0.14
R8106 IREF.n1157 IREF.n789 0.14
R8107 IREF.n1159 IREF.n1158 0.14
R8108 IREF.n1159 IREF.n786 0.14
R8109 IREF.n1184 IREF.n787 0.14
R8110 IREF.n1179 IREF.n787 0.14
R8111 IREF.n1178 IREF.n1177 0.14
R8112 IREF.n1177 IREF.n1167 0.14
R8113 IREF.n1172 IREF.n1171 0.14
R8114 IREF.n1357 IREF.n1349 0.14
R8115 IREF.n1358 IREF.n1357 0.14
R8116 IREF.n1359 IREF.n1347 0.14
R8117 IREF.n1363 IREF.n1347 0.14
R8118 IREF.n1375 IREF.n1368 0.14
R8119 IREF.n1375 IREF.n1374 0.14
R8120 IREF.n5 IREF.n4 0.14
R8121 IREF.n9 IREF.n4 0.14
R8122 IREF.n10 IREF.n3 0.14
R8123 IREF.n13 IREF.n3 0.14
R8124 IREF.n14 IREF.n2 0.14
R8125 IREF.n17 IREF.n2 0.14
R8126 IREF.n1386 IREF.n18 0.14
R8127 IREF.n28 IREF.n27 0.1355
R8128 IREF.n1385 IREF.n19 0.1355
R8129 IREF.n1382 IREF.n1346 0.120905
R8130 IREF.n929 IREF.n928 0.118921
R8131 IREF.n884 IREF.n865 0.118921
R8132 IREF.n1076 IREF.n1054 0.118921
R8133 IREF.n1036 IREF.n1035 0.118921
R8134 IREF.n948 IREF.n947 0.116553
R8135 IREF.n888 IREF.n864 0.116553
R8136 IREF.n1072 IREF.n1055 0.116553
R8137 IREF.n1113 IREF.n1112 0.116553
R8138 IREF.n935 IREF.n933 0.114184
R8139 IREF.n915 IREF.n914 0.114184
R8140 IREF.n894 IREF.n893 0.114184
R8141 IREF.n1067 IREF.n1057 0.114184
R8142 IREF.n1049 IREF.n1047 0.114184
R8143 IREF.n1042 IREF.n1040 0.114184
R8144 IREF.n1244 IREF.n1243 0.109179
R8145 IREF.n1239 IREF.n1238 0.109179
R8146 IREF.n86 IREF.n85 0.109179
R8147 IREF.n92 IREF.n43 0.109179
R8148 IREF.n505 IREF.n504 0.109179
R8149 IREF.n511 IREF.n134 0.109179
R8150 IREF.n436 IREF.n435 0.109179
R8151 IREF.n442 IREF.n392 0.109179
R8152 IREF.n1224 IREF.n1223 0.107155
R8153 IREF.n1258 IREF.n122 0.107155
R8154 IREF.n1280 IREF.n1279 0.107155
R8155 IREF.n70 IREF.n51 0.107155
R8156 IREF.n542 IREF.n541 0.107155
R8157 IREF.n489 IREF.n142 0.107155
R8158 IREF.n461 IREF.n154 0.107155
R8159 IREF.n419 IREF.n418 0.107155
R8160 IREF.n1229 IREF.n1228 0.103632
R8161 IREF.n1261 IREF.n116 0.103632
R8162 IREF.n1285 IREF.n99 0.103632
R8163 IREF.n63 IREF.n62 0.103632
R8164 IREF.n547 IREF.n518 0.103632
R8165 IREF.n482 IREF.n481 0.103632
R8166 IREF.n454 IREF.n453 0.103632
R8167 IREF.n414 IREF.n404 0.103632
R8168 IREF.n321 IREF.n320 0.102991
R8169 IREF.n316 IREF.n315 0.102991
R8170 IREF.n215 IREF.n214 0.102991
R8171 IREF.n221 IREF.n164 0.102991
R8172 IREF.n727 IREF.n726 0.102991
R8173 IREF.n733 IREF.n558 0.102991
R8174 IREF.n646 IREF.n645 0.102991
R8175 IREF.n641 IREF.n640 0.102991
R8176 IREF.n939 IREF.n936 0.0987895
R8177 IREF.n921 IREF.n920 0.0987895
R8178 IREF.n900 IREF.n899 0.0987895
R8179 IREF.n875 IREF.n874 0.0987895
R8180 IREF.n1062 IREF.n1059 0.0987895
R8181 IREF.n1085 IREF.n1050 0.0987895
R8182 IREF.n1104 IREF.n1043 0.0987895
R8183 IREF.n1028 IREF.n1027 0.0987895
R8184 IREF.n305 IREF.n269 0.0933826
R8185 IREF.n350 IREF.n349 0.0933826
R8186 IREF.n379 IREF.n227 0.0933826
R8187 IREF.n185 IREF.n184 0.0933826
R8188 IREF.n774 IREF.n739 0.0933826
R8189 IREF.n697 IREF.n696 0.0933826
R8190 IREF.n662 IREF.n586 0.0933826
R8191 IREF.n609 IREF.n601 0.0933826
R8192 IREF.n297 IREF.n274 0.092742
R8193 IREF.n341 IREF.n340 0.092742
R8194 IREF.n371 IREF.n232 0.092742
R8195 IREF.n194 IREF.n193 0.092742
R8196 IREF.n766 IREF.n744 0.092742
R8197 IREF.n706 IREF.n705 0.092742
R8198 IREF.n671 IREF.n582 0.092742
R8199 IREF.n618 IREF.n597 0.092742
R8200 IREF IREF.n1387 0.0822105
R8201 IREF.n1219 IREF.n1218 0.0821726
R8202 IREF.n1253 IREF.n1252 0.0821726
R8203 IREF.n1275 IREF.n1274 0.0821726
R8204 IREF.n75 IREF.n47 0.0821726
R8205 IREF.n289 IREF.n279 0.0821726
R8206 IREF.n332 IREF.n331 0.0821726
R8207 IREF.n239 IREF.n237 0.0821726
R8208 IREF.n204 IREF.n170 0.0821726
R8209 IREF.n537 IREF.n536 0.0821726
R8210 IREF.n494 IREF.n138 0.0821726
R8211 IREF.n466 IREF.n150 0.0821726
R8212 IREF.n427 IREF.n398 0.0821726
R8213 IREF.n751 IREF.n749 0.0821726
R8214 IREF.n716 IREF.n564 0.0821726
R8215 IREF.n678 IREF.n578 0.0821726
R8216 IREF.n625 IREF.n593 0.0821726
R8217 IREF.n28 IREF.n24 0.0733942
R8218 IREF.n922 IREF.n921 0.0490526
R8219 IREF.n901 IREF.n900 0.0490526
R8220 IREF.n874 IREF.n867 0.0490526
R8221 IREF.n1082 IREF.n1050 0.0490526
R8222 IREF.n1101 IREF.n1043 0.0490526
R8223 IREF.n1029 IREF.n1028 0.0490526
R8224 IREF.n1243 IREF.n1193 0.0426132
R8225 IREF.n1238 IREF.n1237 0.0426132
R8226 IREF.n88 IREF.n86 0.0426132
R8227 IREF.n93 IREF.n92 0.0426132
R8228 IREF.n507 IREF.n505 0.0426132
R8229 IREF.n512 IREF.n511 0.0426132
R8230 IREF.n438 IREF.n436 0.0426132
R8231 IREF.n443 IREF.n442 0.0426132
R8232 IREF.n1245 IREF.n1244 0.0412547
R8233 IREF.n1239 IREF.n1195 0.0412547
R8234 IREF.n85 IREF.n45 0.0412547
R8235 IREF.n87 IREF.n43 0.0412547
R8236 IREF.n504 IREF.n136 0.0412547
R8237 IREF.n506 IREF.n134 0.0412547
R8238 IREF.n435 IREF.n394 0.0412547
R8239 IREF.n437 IREF.n392 0.0412547
R8240 IREF.n1230 IREF.n1229 0.0402153
R8241 IREF.n1225 IREF.n1224 0.0402153
R8242 IREF.n1220 IREF.n1219 0.0402153
R8243 IREF.n1218 IREF.n1212 0.0402153
R8244 IREF.n1265 IREF.n116 0.0402153
R8245 IREF.n1259 IREF.n1258 0.0402153
R8246 IREF.n1254 IREF.n1253 0.0402153
R8247 IREF.n1252 IREF.n129 0.0402153
R8248 IREF.n1286 IREF.n1285 0.0402153
R8249 IREF.n1281 IREF.n1280 0.0402153
R8250 IREF.n1276 IREF.n1275 0.0402153
R8251 IREF.n1274 IREF.n111 0.0402153
R8252 IREF.n62 IREF.n56 0.0402153
R8253 IREF.n66 IREF.n51 0.0402153
R8254 IREF.n75 IREF.n49 0.0402153
R8255 IREF.n79 IREF.n47 0.0402153
R8256 IREF.n320 IREF.n260 0.0402153
R8257 IREF.n315 IREF.n314 0.0402153
R8258 IREF.n217 IREF.n215 0.0402153
R8259 IREF.n222 IREF.n221 0.0402153
R8260 IREF.n548 IREF.n547 0.0402153
R8261 IREF.n543 IREF.n542 0.0402153
R8262 IREF.n538 IREF.n537 0.0402153
R8263 IREF.n536 IREF.n530 0.0402153
R8264 IREF.n481 IREF.n147 0.0402153
R8265 IREF.n485 IREF.n142 0.0402153
R8266 IREF.n494 IREF.n140 0.0402153
R8267 IREF.n498 IREF.n138 0.0402153
R8268 IREF.n453 IREF.n159 0.0402153
R8269 IREF.n457 IREF.n154 0.0402153
R8270 IREF.n466 IREF.n152 0.0402153
R8271 IREF.n470 IREF.n150 0.0402153
R8272 IREF.n409 IREF.n404 0.0402153
R8273 IREF.n418 IREF.n402 0.0402153
R8274 IREF.n423 IREF.n398 0.0402153
R8275 IREF.n428 IREF.n427 0.0402153
R8276 IREF.n729 IREF.n727 0.0402153
R8277 IREF.n734 IREF.n733 0.0402153
R8278 IREF.n645 IREF.n634 0.0402153
R8279 IREF.n640 IREF.n639 0.0402153
R8280 IREF.n322 IREF.n321 0.0389342
R8281 IREF.n316 IREF.n262 0.0389342
R8282 IREF.n214 IREF.n166 0.0389342
R8283 IREF.n216 IREF.n164 0.0389342
R8284 IREF.n726 IREF.n560 0.0389342
R8285 IREF.n728 IREF.n558 0.0389342
R8286 IREF.n647 IREF.n646 0.0389342
R8287 IREF.n641 IREF.n636 0.0389342
R8288 IREF.n285 IREF.n281 0.0338096
R8289 IREF.n330 IREF.n256 0.0338096
R8290 IREF.n363 IREF.n362 0.0338096
R8291 IREF.n205 IREF.n168 0.0338096
R8292 IREF.n758 IREF.n757 0.0338096
R8293 IREF.n717 IREF.n562 0.0338096
R8294 IREF.n684 IREF.n682 0.0338096
R8295 IREF.n631 IREF.n629 0.0338096
R8296 IREF.n941 IREF.n935 0.0336579
R8297 IREF.n916 IREF.n915 0.0336579
R8298 IREF.n893 IREF.n862 0.0336579
R8299 IREF.n872 IREF.n869 0.0336579
R8300 IREF.n1064 IREF.n1057 0.0336579
R8301 IREF.n1087 IREF.n1049 0.0336579
R8302 IREF.n1106 IREF.n1042 0.0336579
R8303 IREF.n1023 IREF.n1022 0.0336579
R8304 IREF.n1215 IREF.n1213 0.0325285
R8305 IREF.n1248 IREF.n1190 0.0325285
R8306 IREF.n1270 IREF.n113 0.0325285
R8307 IREF.n81 IREF.n80 0.0325285
R8308 IREF.n282 IREF.n280 0.0325285
R8309 IREF.n326 IREF.n325 0.0325285
R8310 IREF.n359 IREF.n243 0.0325285
R8311 IREF.n210 IREF.n209 0.0325285
R8312 IREF.n533 IREF.n531 0.0325285
R8313 IREF.n500 IREF.n499 0.0325285
R8314 IREF.n472 IREF.n471 0.0325285
R8315 IREF.n431 IREF.n396 0.0325285
R8316 IREF.n755 IREF.n754 0.0325285
R8317 IREF.n722 IREF.n721 0.0325285
R8318 IREF.n687 IREF.n576 0.0325285
R8319 IREF.n650 IREF.n591 0.0325285
R8320 IREF.n1233 IREF.n1198 0.0318879
R8321 IREF.n1267 IREF.n1266 0.0318879
R8322 IREF.n1288 IREF.n1287 0.0318879
R8323 IREF.n59 IREF.n58 0.0318879
R8324 IREF.n550 IREF.n549 0.0318879
R8325 IREF.n477 IREF.n476 0.0318879
R8326 IREF.n449 IREF.n448 0.0318879
R8327 IREF.n407 IREF.n406 0.0318879
R8328 IREF.n947 IREF.n946 0.0312895
R8329 IREF.n909 IREF.n858 0.0312895
R8330 IREF.n891 IREF.n864 0.0312895
R8331 IREF.n1069 IREF.n1055 0.0312895
R8332 IREF.n1093 IREF.n1092 0.0312895
R8333 IREF.n1112 IREF.n1111 0.0312895
R8334 IREF.n1228 IREF.n1202 0.0312473
R8335 IREF.n1261 IREF.n1260 0.0312473
R8336 IREF.n101 IREF.n99 0.0312473
R8337 IREF.n63 IREF.n54 0.0312473
R8338 IREF.n520 IREF.n518 0.0312473
R8339 IREF.n482 IREF.n145 0.0312473
R8340 IREF.n454 IREF.n157 0.0312473
R8341 IREF.n414 IREF.n405 0.0312473
R8342 IREF.n310 IREF.n309 0.0306068
R8343 IREF.n306 IREF.n268 0.0306068
R8344 IREF.n356 IREF.n355 0.0306068
R8345 IREF.n353 IREF.n245 0.0306068
R8346 IREF.n386 IREF.n162 0.0306068
R8347 IREF.n383 IREF.n382 0.0306068
R8348 IREF.n181 IREF.n178 0.0306068
R8349 IREF.n781 IREF.n556 0.0306068
R8350 IREF.n778 IREF.n777 0.0306068
R8351 IREF.n691 IREF.n574 0.0306068
R8352 IREF.n693 IREF.n572 0.0306068
R8353 IREF.n655 IREF.n654 0.0306068
R8354 IREF.n659 IREF.n658 0.0306068
R8355 IREF.n606 IREF.n605 0.0306068
R8356 IREF.n302 IREF.n301 0.0299662
R8357 IREF.n298 IREF.n273 0.0299662
R8358 IREF.n346 IREF.n247 0.0299662
R8359 IREF.n344 IREF.n250 0.0299662
R8360 IREF.n378 IREF.n229 0.0299662
R8361 IREF.n375 IREF.n374 0.0299662
R8362 IREF.n188 IREF.n176 0.0299662
R8363 IREF.n190 IREF.n174 0.0299662
R8364 IREF.n773 IREF.n741 0.0299662
R8365 IREF.n770 IREF.n769 0.0299662
R8366 IREF.n700 IREF.n570 0.0299662
R8367 IREF.n702 IREF.n568 0.0299662
R8368 IREF.n664 IREF.n663 0.0299662
R8369 IREF.n668 IREF.n667 0.0299662
R8370 IREF.n611 IREF.n610 0.0299662
R8371 IREF.n615 IREF.n614 0.0299662
R8372 IREF.n928 IREF.n927 0.0289211
R8373 IREF.n907 IREF.n906 0.0289211
R8374 IREF.n881 IREF.n865 0.0289211
R8375 IREF.n1054 IREF.n1052 0.0289211
R8376 IREF.n1095 IREF.n1045 0.0289211
R8377 IREF.n1035 IREF.n1034 0.0289211
R8378 IREF.n1223 IREF.n1207 0.0270836
R8379 IREF.n124 IREF.n122 0.0270836
R8380 IREF.n1279 IREF.n106 0.0270836
R8381 IREF.n70 IREF.n52 0.0270836
R8382 IREF.n541 IREF.n525 0.0270836
R8383 IREF.n489 IREF.n143 0.0270836
R8384 IREF.n461 IREF.n155 0.0270836
R8385 IREF.n419 IREF.n400 0.0270836
R8386 IREF.n294 IREF.n293 0.0258025
R8387 IREF.n290 IREF.n278 0.0258025
R8388 IREF.n337 IREF.n252 0.0258025
R8389 IREF.n335 IREF.n254 0.0258025
R8390 IREF.n370 IREF.n234 0.0258025
R8391 IREF.n367 IREF.n366 0.0258025
R8392 IREF.n197 IREF.n172 0.0258025
R8393 IREF.n200 IREF.n199 0.0258025
R8394 IREF.n765 IREF.n746 0.0258025
R8395 IREF.n762 IREF.n761 0.0258025
R8396 IREF.n709 IREF.n566 0.0258025
R8397 IREF.n712 IREF.n711 0.0258025
R8398 IREF.n674 IREF.n673 0.0258025
R8399 IREF.n679 IREF.n580 0.0258025
R8400 IREF.n621 IREF.n620 0.0258025
R8401 IREF.n626 IREF.n595 0.0258025
R8402 IREF.n180 IREF.n179 0.0170406
R8403 IREF.n603 IREF.n602 0.0170406
R8404 IREF.n294 IREF.n274 0.0149128
R8405 IREF.n290 IREF.n289 0.0149128
R8406 IREF.n340 IREF.n252 0.0149128
R8407 IREF.n332 IREF.n254 0.0149128
R8408 IREF.n371 IREF.n370 0.0149128
R8409 IREF.n366 IREF.n237 0.0149128
R8410 IREF.n194 IREF.n172 0.0149128
R8411 IREF.n199 IREF.n170 0.0149128
R8412 IREF.n766 IREF.n765 0.0149128
R8413 IREF.n761 IREF.n749 0.0149128
R8414 IREF.n706 IREF.n566 0.0149128
R8415 IREF.n711 IREF.n564 0.0149128
R8416 IREF.n674 IREF.n671 0.0149128
R8417 IREF.n679 IREF.n678 0.0149128
R8418 IREF.n621 IREF.n618 0.0149128
R8419 IREF.n626 IREF.n625 0.0149128
R8420 IREF.n1220 IREF.n1207 0.0136317
R8421 IREF.n1254 IREF.n124 0.0136317
R8422 IREF.n1276 IREF.n106 0.0136317
R8423 IREF.n52 IREF.n49 0.0136317
R8424 IREF.n278 IREF.n276 0.0136317
R8425 IREF.n336 IREF.n335 0.0136317
R8426 IREF.n367 IREF.n236 0.0136317
R8427 IREF.n200 IREF.n198 0.0136317
R8428 IREF.n538 IREF.n525 0.0136317
R8429 IREF.n143 IREF.n140 0.0136317
R8430 IREF.n155 IREF.n152 0.0136317
R8431 IREF.n423 IREF.n400 0.0136317
R8432 IREF.n762 IREF.n748 0.0136317
R8433 IREF.n712 IREF.n710 0.0136317
R8434 IREF.n672 IREF.n580 0.0136317
R8435 IREF.n619 IREF.n595 0.0136317
R8436 IREF.n302 IREF.n269 0.0107491
R8437 IREF.n298 IREF.n297 0.0107491
R8438 IREF.n349 IREF.n247 0.0107491
R8439 IREF.n341 IREF.n250 0.0107491
R8440 IREF.n379 IREF.n378 0.0107491
R8441 IREF.n374 IREF.n232 0.0107491
R8442 IREF.n185 IREF.n176 0.0107491
R8443 IREF.n193 IREF.n174 0.0107491
R8444 IREF.n774 IREF.n773 0.0107491
R8445 IREF.n769 IREF.n744 0.0107491
R8446 IREF.n697 IREF.n570 0.0107491
R8447 IREF.n705 IREF.n568 0.0107491
R8448 IREF.n664 IREF.n662 0.0107491
R8449 IREF.n668 IREF.n582 0.0107491
R8450 IREF.n611 IREF.n609 0.0107491
R8451 IREF.n615 IREF.n597 0.0107491
R8452 IREF.n306 IREF.n305 0.0101085
R8453 IREF.n350 IREF.n245 0.0101085
R8454 IREF.n382 IREF.n227 0.0101085
R8455 IREF.n184 IREF.n178 0.0101085
R8456 IREF.n777 IREF.n739 0.0101085
R8457 IREF.n696 IREF.n572 0.0101085
R8458 IREF.n659 IREF.n586 0.0101085
R8459 IREF.n606 IREF.n601 0.0101085
R8460 IREF.n1225 IREF.n1202 0.00946797
R8461 IREF.n1260 IREF.n1259 0.00946797
R8462 IREF.n1281 IREF.n101 0.00946797
R8463 IREF.n66 IREF.n54 0.00946797
R8464 IREF.n273 IREF.n271 0.00946797
R8465 IREF.n345 IREF.n344 0.00946797
R8466 IREF.n375 IREF.n231 0.00946797
R8467 IREF.n190 IREF.n189 0.00946797
R8468 IREF.n543 IREF.n520 0.00946797
R8469 IREF.n485 IREF.n145 0.00946797
R8470 IREF.n457 IREF.n157 0.00946797
R8471 IREF.n405 IREF.n402 0.00946797
R8472 IREF.n770 IREF.n743 0.00946797
R8473 IREF.n702 IREF.n701 0.00946797
R8474 IREF.n667 IREF.n584 0.00946797
R8475 IREF.n614 IREF.n599 0.00946797
R8476 IREF.n1230 IREF.n1198 0.0088274
R8477 IREF.n1266 IREF.n1265 0.0088274
R8478 IREF.n1287 IREF.n1286 0.0088274
R8479 IREF.n58 IREF.n56 0.0088274
R8480 IREF.n268 IREF.n266 0.0088274
R8481 IREF.n354 IREF.n353 0.0088274
R8482 IREF.n383 IREF.n226 0.0088274
R8483 IREF.n181 IREF.n180 0.0088274
R8484 IREF.n549 IREF.n548 0.0088274
R8485 IREF.n476 IREF.n147 0.0088274
R8486 IREF.n448 IREF.n159 0.0088274
R8487 IREF.n409 IREF.n407 0.0088274
R8488 IREF.n778 IREF.n738 0.0088274
R8489 IREF.n693 IREF.n692 0.0088274
R8490 IREF.n658 IREF.n588 0.0088274
R8491 IREF.n605 IREF.n603 0.0088274
R8492 IREF.n1213 IREF.n1212 0.00818683
R8493 IREF.n1190 IREF.n129 0.00818683
R8494 IREF.n113 IREF.n111 0.00818683
R8495 IREF.n80 IREF.n79 0.00818683
R8496 IREF.n531 IREF.n530 0.00818683
R8497 IREF.n499 IREF.n498 0.00818683
R8498 IREF.n471 IREF.n470 0.00818683
R8499 IREF.n428 IREF.n396 0.00818683
R8500 IREF.n281 IREF.n279 0.00690569
R8501 IREF.n285 IREF.n284 0.00690569
R8502 IREF.n331 IREF.n330 0.00690569
R8503 IREF.n327 IREF.n256 0.00690569
R8504 IREF.n363 IREF.n239 0.00690569
R8505 IREF.n362 IREF.n240 0.00690569
R8506 IREF.n205 IREF.n204 0.00690569
R8507 IREF.n208 IREF.n168 0.00690569
R8508 IREF.n758 IREF.n751 0.00690569
R8509 IREF.n757 IREF.n752 0.00690569
R8510 IREF.n717 IREF.n716 0.00690569
R8511 IREF.n720 IREF.n562 0.00690569
R8512 IREF.n682 IREF.n578 0.00690569
R8513 IREF.n684 IREF.n683 0.00690569
R8514 IREF.n629 IREF.n593 0.00690569
R8515 IREF.n631 IREF.n630 0.00690569
R8516 IREF.n1182 IREF.n1181 0.00523684
R8517 IREF.n1176 IREF.n1175 0.00523684
R8518 IREF.n1169 IREF.n1168 0.00523684
R8519 IREF.n1149 IREF.n1148 0.00523684
R8520 IREF.n1155 IREF.n1154 0.00523684
R8521 IREF.n1161 IREF.n1160 0.00523684
R8522 IREF.n1125 IREF.n798 0.00523684
R8523 IREF.n1130 IREF.n796 0.00523684
R8524 IREF.n1136 IREF.n1135 0.00523684
R8525 IREF.n1142 IREF.n1141 0.00523684
R8526 IREF.n809 IREF.n802 0.00523684
R8527 IREF.n814 IREF.n800 0.00523684
R8528 IREF.n955 IREF.n953 0.00523684
R8529 IREF.n966 IREF.n956 0.00523684
R8530 IREF.n961 IREF.n958 0.00523684
R8531 IREF.n848 IREF.n846 0.00523684
R8532 IREF.n984 IREF.n849 0.00523684
R8533 IREF.n979 IREF.n851 0.00523684
R8534 IREF.n1011 IREF.n1010 0.00523684
R8535 IREF.n1005 IREF.n1004 0.00523684
R8536 IREF.n843 IREF.n841 0.00523684
R8537 IREF.n996 IREF.n844 0.00523684
R8538 IREF.n828 IREF.n827 0.00523684
R8539 IREF.n834 IREF.n833 0.00523684
R8540 IREF.n1356 IREF.n1355 0.00523684
R8541 IREF.n1362 IREF.n1361 0.00523684
R8542 IREF.n1386 IREF.n1385 0.005
R8543 IREF.n1195 IREF.n1193 0.00185849
R8544 IREF.n1237 IREF.n1196 0.00185849
R8545 IREF.n88 IREF.n87 0.00185849
R8546 IREF.n94 IREF.n93 0.00185849
R8547 IREF.n507 IREF.n506 0.00185849
R8548 IREF.n513 IREF.n512 0.00185849
R8549 IREF.n438 IREF.n437 0.00185849
R8550 IREF.n444 IREF.n443 0.00185849
R8551 IREF.n309 IREF.n266 0.00178114
R8552 IREF.n301 IREF.n271 0.00178114
R8553 IREF.n293 IREF.n276 0.00178114
R8554 IREF.n284 IREF.n282 0.00178114
R8555 IREF.n355 IREF.n354 0.00178114
R8556 IREF.n346 IREF.n345 0.00178114
R8557 IREF.n337 IREF.n336 0.00178114
R8558 IREF.n327 IREF.n326 0.00178114
R8559 IREF.n226 IREF.n162 0.00178114
R8560 IREF.n231 IREF.n229 0.00178114
R8561 IREF.n236 IREF.n234 0.00178114
R8562 IREF.n243 IREF.n240 0.00178114
R8563 IREF.n262 IREF.n260 0.00178114
R8564 IREF.n314 IREF.n263 0.00178114
R8565 IREF.n217 IREF.n216 0.00178114
R8566 IREF.n223 IREF.n222 0.00178114
R8567 IREF.n189 IREF.n188 0.00178114
R8568 IREF.n198 IREF.n197 0.00178114
R8569 IREF.n209 IREF.n208 0.00178114
R8570 IREF.n738 IREF.n556 0.00178114
R8571 IREF.n743 IREF.n741 0.00178114
R8572 IREF.n748 IREF.n746 0.00178114
R8573 IREF.n754 IREF.n752 0.00178114
R8574 IREF.n692 IREF.n691 0.00178114
R8575 IREF.n701 IREF.n700 0.00178114
R8576 IREF.n710 IREF.n709 0.00178114
R8577 IREF.n721 IREF.n720 0.00178114
R8578 IREF.n654 IREF.n588 0.00178114
R8579 IREF.n663 IREF.n584 0.00178114
R8580 IREF.n673 IREF.n672 0.00178114
R8581 IREF.n683 IREF.n576 0.00178114
R8582 IREF.n729 IREF.n728 0.00178114
R8583 IREF.n735 IREF.n734 0.00178114
R8584 IREF.n636 IREF.n634 0.00178114
R8585 IREF.n639 IREF.n637 0.00178114
R8586 IREF.n610 IREF.n599 0.00178114
R8587 IREF.n620 IREF.n619 0.00178114
R8588 IREF.n630 IREF.n591 0.00178114
R8589 IREF.n35 IREF.n34 0.00168421
R8590 IREF.n16 IREF.n15 0.00168421
R8591 IREF.n12 IREF.n11 0.00168421
R8592 IREF.n8 IREF.n7 0.00168421
R8593 IREF.n1387 IREF.n1 0.00168421
R8594 a_n11737_n15980.n130 a_n11737_n15980.n129 12.734
R8595 a_n11737_n15980.n56 a_n11737_n15980.t27 8.41809
R8596 a_n11737_n15980.n57 a_n11737_n15980.t36 8.41809
R8597 a_n11737_n15980.n56 a_n11737_n15980.t44 8.37125
R8598 a_n11737_n15980.n60 a_n11737_n15980.t63 8.37125
R8599 a_n11737_n15980.n57 a_n11737_n15980.t48 8.37125
R8600 a_n11737_n15980.n103 a_n11737_n15980.t29 8.33806
R8601 a_n11737_n15980.n97 a_n11737_n15980.t62 8.3366
R8602 a_n11737_n15980.n82 a_n11737_n15980.t56 8.26493
R8603 a_n11737_n15980.n116 a_n11737_n15980.t39 8.2602
R8604 a_n11737_n15980.n17 a_n11737_n15980.t35 8.06917
R8605 a_n11737_n15980.n28 a_n11737_n15980.t42 8.06917
R8606 a_n11737_n15980.n13 a_n11737_n15980.t28 8.06917
R8607 a_n11737_n15980.n13 a_n11737_n15980.t41 8.06917
R8608 a_n11737_n15980.n11 a_n11737_n15980.t53 8.06917
R8609 a_n11737_n15980.n11 a_n11737_n15980.t40 8.06917
R8610 a_n11737_n15980.n62 a_n11737_n15980.t52 8.06917
R8611 a_n11737_n15980.n17 a_n11737_n15980.t64 8.06917
R8612 a_n11737_n15980.n30 a_n11737_n15980.t34 8.06917
R8613 a_n11737_n15980.n7 a_n11737_n15980.t50 8.06917
R8614 a_n11737_n15980.n7 a_n11737_n15980.t37 8.06917
R8615 a_n11737_n15980.n32 a_n11737_n15980.t49 8.06917
R8616 a_n11737_n15980.n76 a_n11737_n15980.t55 8.06917
R8617 a_n11737_n15980.n3 a_n11737_n15980.t45 8.06917
R8618 a_n11737_n15980.n3 a_n11737_n15980.t54 8.06917
R8619 a_n11737_n15980.n21 a_n11737_n15980.t26 8.06917
R8620 a_n11737_n15980.n21 a_n11737_n15980.t58 8.06917
R8621 a_n11737_n15980.n70 a_n11737_n15980.t25 8.06917
R8622 a_n11737_n15980.n96 a_n11737_n15980.t51 8.06917
R8623 a_n11737_n15980.n0 a_n11737_n15980.t61 8.06917
R8624 a_n11737_n15980.n94 a_n11737_n15980.t32 8.06917
R8625 a_n11737_n15980.n93 a_n11737_n15980.t60 8.06917
R8626 a_n11737_n15980.n92 a_n11737_n15980.t31 8.06917
R8627 a_n11737_n15980.n90 a_n11737_n15980.t57 8.06917
R8628 a_n11737_n15980.n83 a_n11737_n15980.t43 8.06917
R8629 a_n11737_n15980.n110 a_n11737_n15980.t30 8.06917
R8630 a_n11737_n15980.n104 a_n11737_n15980.t59 8.06917
R8631 a_n11737_n15980.n112 a_n11737_n15980.t46 8.06917
R8632 a_n11737_n15980.n113 a_n11737_n15980.t33 8.06917
R8633 a_n11737_n15980.n114 a_n11737_n15980.t47 8.06917
R8634 a_n11737_n15980.n117 a_n11737_n15980.t24 8.06917
R8635 a_n11737_n15980.n123 a_n11737_n15980.t38 8.06917
R8636 a_n11737_n15980.n59 a_n11737_n15980.t0 6.65728
R8637 a_n11737_n15980.n45 a_n11737_n15980.t13 6.51495
R8638 a_n11737_n15980.n133 a_n11737_n15980.t11 6.40828
R8639 a_n11737_n15980.n42 a_n11737_n15980.t22 6.37877
R8640 a_n11737_n15980.n59 a_n11737_n15980.t1 5.74368
R8641 a_n11737_n15980.n46 a_n11737_n15980.t15 5.24318
R8642 a_n11737_n15980.n64 a_n11737_n15980.n31 2.4223
R8643 a_n11737_n15980.n71 a_n11737_n15980.n33 2.42484
R8644 a_n11737_n15980.n72 a_n11737_n15980.n33 2.4256
R8645 a_n11737_n15980.n39 a_n11737_n15980.n38 2.24636
R8646 a_n11737_n15980.t12 a_n11737_n15980.n35 5.26436
R8647 a_n11737_n15980.n53 a_n11737_n15980.n42 4.60825
R8648 a_n11737_n15980.n34 a_n11737_n15980.n141 3.79435
R8649 a_n11737_n15980.n38 a_n11737_n15980.n133 4.59811
R8650 a_n11737_n15980.n22 a_n11737_n15980.n21 0.592766
R8651 a_n11737_n15980.n12 a_n11737_n15980.n11 0.592803
R8652 a_n11737_n15980.n15 a_n11737_n15980.n13 0.591918
R8653 a_n11737_n15980.n17 a_n11737_n15980.n18 0.591826
R8654 a_n11737_n15980.n37 a_n11737_n15980.n36 2.24389
R8655 a_n11737_n15980.n49 a_n11737_n15980.n43 4.5005
R8656 a_n11737_n15980.n10 a_n11737_n15980.n66 4.5005
R8657 a_n11737_n15980.n13 a_n11737_n15980.n14 0.591264
R8658 a_n11737_n15980.n67 a_n11737_n15980.n24 4.5005
R8659 a_n11737_n15980.n31 a_n11737_n15980.n30 0.0133501
R8660 a_n11737_n15980.n16 a_n11737_n15980.n64 4.5005
R8661 a_n11737_n15980.n19 a_n11737_n15980.n17 0.604195
R8662 a_n11737_n15980.n29 a_n11737_n15980.n63 4.5005
R8663 a_n11737_n15980.n69 a_n11737_n15980.n68 4.5005
R8664 a_n11737_n15980.n28 a_n11737_n15980.n27 0.0143905
R8665 a_n11737_n15980.n20 a_n11737_n15980.n74 4.5005
R8666 a_n11737_n15980.n2 a_n11737_n15980.n75 4.5005
R8667 a_n11737_n15980.n3 a_n11737_n15980.n4 0.591675
R8668 a_n11737_n15980.n9 a_n11737_n15980.n7 0.604671
R8669 a_n11737_n15980.n6 a_n11737_n15980.n71 4.5005
R8670 a_n11737_n15980.n32 a_n11737_n15980.n33 0.0107891
R8671 a_n11737_n15980.n7 a_n11737_n15980.n8 0.604671
R8672 a_n11737_n15980.n72 a_n11737_n15980.n6 4.5005
R8673 a_n11737_n15980.n2 a_n11737_n15980.n23 4.5005
R8674 a_n11737_n15980.n5 a_n11737_n15980.n3 0.591675
R8675 a_n11737_n15980.n84 a_n11737_n15980.n81 4.5005
R8676 a_n11737_n15980.n86 a_n11737_n15980.n85 4.5005
R8677 a_n11737_n15980.n87 a_n11737_n15980.n80 4.5005
R8678 a_n11737_n15980.n89 a_n11737_n15980.n88 4.5005
R8679 a_n11737_n15980.n91 a_n11737_n15980.n79 4.5005
R8680 a_n11737_n15980.n1 a_n11737_n15980.n0 1.44113
R8681 a_n11737_n15980.n98 a_n11737_n15980.n95 4.5005
R8682 a_n11737_n15980.n111 a_n11737_n15980.n100 4.5005
R8683 a_n11737_n15980.n109 a_n11737_n15980.n108 4.5005
R8684 a_n11737_n15980.n107 a_n11737_n15980.n102 4.5005
R8685 a_n11737_n15980.n106 a_n11737_n15980.n105 4.5005
R8686 a_n11737_n15980.n126 a_n11737_n15980.n125 4.5005
R8687 a_n11737_n15980.n124 a_n11737_n15980.n101 4.5005
R8688 a_n11737_n15980.n122 a_n11737_n15980.n121 4.5005
R8689 a_n11737_n15980.n120 a_n11737_n15980.n115 4.5005
R8690 a_n11737_n15980.n119 a_n11737_n15980.n118 4.5005
R8691 a_n11737_n15980.n140 a_n11737_n15980.n139 4.5005
R8692 a_n11737_n15980.n40 a_n11737_n15980.n41 2.23676
R8693 a_n11737_n15980.n36 a_n11737_n15980.t7 3.79594
R8694 a_n11737_n15980.t23 a_n11737_n15980.n40 3.79475
R8695 a_n11737_n15980.n138 a_n11737_n15980.t19 3.77936
R8696 a_n11737_n15980.n50 a_n11737_n15980.t5 3.77818
R8697 a_n11737_n15980.n45 a_n11737_n15980.n44 3.77318
R8698 a_n11737_n15980.n136 a_n11737_n15980.n135 3.77081
R8699 a_n11737_n15980.n48 a_n11737_n15980.n47 3.75571
R8700 a_n11737_n15980.n131 a_n11737_n15980.n55 2.69513
R8701 a_n11737_n15980.n77 a_n11737_n15980.n75 2.4256
R8702 a_n11737_n15980.n23 a_n11737_n15980.n77 2.42484
R8703 a_n11737_n15980.n31 a_n11737_n15980.n63 2.43326
R8704 a_n11737_n15980.n38 a_n11737_n15980.n134 2.32949
R8705 a_n11737_n15980.n128 a_n11737_n15980.n99 2.30989
R8706 a_n11737_n15980.n53 a_n11737_n15980.n52 2.30818
R8707 a_n11737_n15980.n138 a_n11737_n15980.n137 2.24481
R8708 a_n11737_n15980.n54 a_n11737_n15980.n53 2.2442
R8709 a_n11737_n15980.n51 a_n11737_n15980.n50 2.24358
R8710 a_n11737_n15980.n73 a_n11737_n15980.n70 2.23529
R8711 a_n11737_n15980.n65 a_n11737_n15980.n62 2.23423
R8712 a_n11737_n15980.n99 a_n11737_n15980.n79 2.18975
R8713 a_n11737_n15980.n127 a_n11737_n15980.n100 2.16725
R8714 a_n11737_n15980.n26 a_n11737_n15980.n5 2.4981
R8715 a_n11737_n15980.n129 a_n11737_n15980.n78 2.07557
R8716 a_n11737_n15980.n78 a_n11737_n15980.n25 2.07182
R8717 a_n11737_n15980.n25 a_n11737_n15980.n15 2.4644
R8718 a_n11737_n15980.n60 a_n11737_n15980.n59 1.7613
R8719 a_n11737_n15980.n58 a_n11737_n15980.n56 1.55888
R8720 a_n11737_n15980.n78 a_n11737_n15980.n26 1.5005
R8721 a_n11737_n15980.n128 a_n11737_n15980.n127 1.5005
R8722 a_n11737_n15980.n58 a_n11737_n15980.n57 1.5005
R8723 a_n11737_n15980.n61 a_n11737_n15980.n60 1.5005
R8724 a_n11737_n15980.n132 a_n11737_n15980.n131 1.5005
R8725 a_n11737_n15980.n141 a_n11737_n15980.t8 1.4705
R8726 a_n11737_n15980.n141 a_n11737_n15980.t14 1.4705
R8727 a_n11737_n15980.n47 a_n11737_n15980.t3 1.4705
R8728 a_n11737_n15980.n47 a_n11737_n15980.t2 1.4705
R8729 a_n11737_n15980.n44 a_n11737_n15980.t18 1.4705
R8730 a_n11737_n15980.n44 a_n11737_n15980.t6 1.4705
R8731 a_n11737_n15980.n52 a_n11737_n15980.t10 1.4705
R8732 a_n11737_n15980.n52 a_n11737_n15980.t9 1.4705
R8733 a_n11737_n15980.n134 a_n11737_n15980.t17 1.4705
R8734 a_n11737_n15980.n134 a_n11737_n15980.t16 1.4705
R8735 a_n11737_n15980.n135 a_n11737_n15980.t4 1.4705
R8736 a_n11737_n15980.n135 a_n11737_n15980.t21 1.4705
R8737 a_n11737_n15980.n82 a_n11737_n15980.n81 1.39514
R8738 a_n11737_n15980.n119 a_n11737_n15980.n116 1.39105
R8739 a_n11737_n15980.n129 a_n11737_n15980.n128 1.35453
R8740 a_n11737_n15980.n46 a_n11737_n15980.n45 1.27228
R8741 a_n11737_n15980.n92 a_n11737_n15980.n91 1.26997
R8742 a_n11737_n15980.n0 a_n11737_n15980.n94 1.24392
R8743 a_n11737_n15980.n112 a_n11737_n15980.n111 1.24204
R8744 a_n11737_n15980.n137 a_n11737_n15980.n136 1.20603
R8745 a_n11737_n15980.n125 a_n11737_n15980.n114 1.20414
R8746 a_n11737_n15980.n98 a_n11737_n15980.n97 1.14132
R8747 a_n11737_n15980.n54 a_n11737_n15980.n51 1.13952
R8748 a_n11737_n15980.n106 a_n11737_n15980.n103 1.13598
R8749 a_n11737_n15980.n37 a_n11737_n15980.n48 1.20574
R8750 a_n11737_n15980.n41 a_n11737_n15980.n34 1.24017
R8751 a_n11737_n15980.n131 a_n11737_n15980.n130 0.963743
R8752 a_n11737_n15980.n48 a_n11737_n15980.n46 0.937067
R8753 a_n11737_n15980.n99 a_n11737_n15980.n1 0.888471
R8754 a_n11737_n15980.n127 a_n11737_n15980.n126 0.71825
R8755 a_n11737_n15980.n93 a_n11737_n15980.n92 0.663658
R8756 a_n11737_n15980.n94 a_n11737_n15980.n93 0.663658
R8757 a_n11737_n15980.n114 a_n11737_n15980.n113 0.655156
R8758 a_n11737_n15980.n113 a_n11737_n15980.n112 0.655156
R8759 a_n11737_n15980.n117 a_n11737_n15980.n116 0.439529
R8760 a_n11737_n15980.n83 a_n11737_n15980.n82 0.432797
R8761 a_n11737_n15980.n122 a_n11737_n15980.n115 0.379447
R8762 a_n11737_n15980.n105 a_n11737_n15980.n102 0.379447
R8763 a_n11737_n15980.n64 a_n11737_n15980.n19 0.745981
R8764 a_n11737_n15980.n9 a_n11737_n15980.n71 0.745252
R8765 a_n11737_n15980.n8 a_n11737_n15980.n72 0.745252
R8766 a_n11737_n15980.n1 a_n11737_n15980.n98 0.498861
R8767 a_n11737_n15980.n66 a_n11737_n15980.n12 0.756573
R8768 a_n11737_n15980.n18 a_n11737_n15980.n63 0.756388
R8769 a_n11737_n15980.n15 a_n11737_n15980.n69 0.756711
R8770 a_n11737_n15980.n74 a_n11737_n15980.n22 0.756011
R8771 a_n11737_n15980.n107 a_n11737_n15980.n106 0.3605
R8772 a_n11737_n15980.n121 a_n11737_n15980.n120 0.3605
R8773 a_n11737_n15980.n97 a_n11737_n15980.n96 0.335806
R8774 a_n11737_n15980.n104 a_n11737_n15980.n103 0.33475
R8775 a_n11737_n15980.n85 a_n11737_n15980.n80 0.302474
R8776 a_n11737_n15980.n87 a_n11737_n15980.n86 0.287375
R8777 a_n11737_n15980.n130 a_n11737_n15980.n61 0.277797
R8778 a_n11737_n15980.n66 a_n11737_n15980.n65 0.208888
R8779 a_n11737_n15980.n74 a_n11737_n15980.n73 0.20887
R8780 a_n11737_n15980.n51 a_n11737_n15980.n43 0.208394
R8781 a_n11737_n15980.n140 a_n11737_n15980.n137 0.208357
R8782 a_n11737_n15980.n61 a_n11737_n15980.n58 0.168946
R8783 a_n11737_n15980.n37 a_n11737_n15980.n43 0.233116
R8784 a_n11737_n15980.n85 a_n11737_n15980.n84 0.147342
R8785 a_n11737_n15980.n89 a_n11737_n15980.n80 0.147342
R8786 a_n11737_n15980.n125 a_n11737_n15980.n124 0.147342
R8787 a_n11737_n15980.n118 a_n11737_n15980.n115 0.147342
R8788 a_n11737_n15980.n109 a_n11737_n15980.n102 0.147342
R8789 a_n11737_n15980.n41 a_n11737_n15980.n140 0.211956
R8790 a_n11737_n15980.n139 a_n11737_n15980.n40 0.142388
R8791 a_n11737_n15980.n55 a_n11737_n15980.n42 0.14
R8792 a_n11737_n15980.n65 a_n11737_n15980.n19 1.12746
R8793 a_n11737_n15980.n14 a_n11737_n15980.n12 1.49123
R8794 a_n11737_n15980.n14 a_n11737_n15980.n24 0.772202
R8795 a_n11737_n15980.n18 a_n11737_n15980.n25 1.21369
R8796 a_n11737_n15980.n69 a_n11737_n15980.n27 2.42126
R8797 a_n11737_n15980.n73 a_n11737_n15980.n9 1.12837
R8798 a_n11737_n15980.n4 a_n11737_n15980.n22 1.49118
R8799 a_n11737_n15980.n75 a_n11737_n15980.n4 0.772883
R8800 a_n11737_n15980.n8 a_n11737_n15980.n26 1.21186
R8801 a_n11737_n15980.n5 a_n11737_n15980.n23 0.772883
R8802 a_n11737_n15980.n86 a_n11737_n15980.n81 0.14
R8803 a_n11737_n15980.n88 a_n11737_n15980.n87 0.14
R8804 a_n11737_n15980.n88 a_n11737_n15980.n79 0.14
R8805 a_n11737_n15980.n108 a_n11737_n15980.n107 0.14
R8806 a_n11737_n15980.n108 a_n11737_n15980.n100 0.14
R8807 a_n11737_n15980.n126 a_n11737_n15980.n101 0.14
R8808 a_n11737_n15980.n121 a_n11737_n15980.n101 0.14
R8809 a_n11737_n15980.n120 a_n11737_n15980.n119 0.14
R8810 a_n11737_n15980.n35 a_n11737_n15980.n39 1.19679
R8811 a_n11737_n15980.n136 a_n11737_n15980.n35 0.932624
R8812 a_n11737_n15980.t20 a_n11737_n15980.n34 6.53226
R8813 a_n11737_n15980.n111 a_n11737_n15980.n110 0.137868
R8814 a_n11737_n15980.n49 a_n11737_n15980.n36 0.137318
R8815 a_n11737_n15980.n133 a_n11737_n15980.n132 0.131
R8816 a_n11737_n15980.n96 a_n11737_n15980.n95 0.128395
R8817 a_n11737_n15980.n105 a_n11737_n15980.n104 0.128395
R8818 a_n11737_n15980.n123 a_n11737_n15980.n122 0.118921
R8819 a_n11737_n15980.n91 a_n11737_n15980.n90 0.114184
R8820 a_n11737_n15980.n50 a_n11737_n15980.n49 0.110782
R8821 a_n11737_n15980.n139 a_n11737_n15980.n138 0.105711
R8822 a_n11737_n15980.n55 a_n11737_n15980.n54 0.0688756
R8823 a_n11737_n15980.n32 a_n11737_n15980.n6 0.0402153
R8824 a_n11737_n15980.n84 a_n11737_n15980.n83 0.0348421
R8825 a_n11737_n15980.n20 a_n11737_n15980.n70 0.0344623
R8826 a_n11737_n15980.n90 a_n11737_n15980.n89 0.0336579
R8827 a_n11737_n15980.n10 a_n11737_n15980.n62 0.0325285
R8828 a_n11737_n15980.n30 a_n11737_n15980.n29 0.0299662
R8829 a_n11737_n15980.n124 a_n11737_n15980.n123 0.0289211
R8830 a_n11737_n15980.n2 a_n11737_n15980.n76 0.0283648
R8831 a_n11737_n15980.n67 a_n11737_n15980.n28 0.0258025
R8832 a_n11737_n15980.n77 a_n11737_n15980.n76 0.0226397
R8833 a_n11737_n15980.n118 a_n11737_n15980.n117 0.0194474
R8834 a_n11737_n15980.n68 a_n11737_n15980.n67 0.0149128
R8835 a_n11737_n15980.n16 a_n11737_n15980.n29 0.0107491
R8836 a_n11737_n15980.n110 a_n11737_n15980.n109 0.00997368
R8837 a_n11737_n15980.n132 a_n11737_n15980.n39 0.0777922
R8838 a_n11737_n15980.n24 a_n11737_n15980.n27 2.43637
R8839 a_n11737_n15980.n0 a_n11737_n15980.n95 0.6755
R8840 a_n11737_n15980.n3 a_n11737_n15980.n2 0.369148
R8841 a_n11737_n15980.n68 a_n11737_n15980.n13 0.354735
R8842 a_n11737_n15980.n7 a_n11737_n15980.n6 0.347689
R8843 a_n11737_n15980.n17 a_n11737_n15980.n16 0.347689
R8844 a_n11737_n15980.n21 a_n11737_n15980.n20 0.346915
R8845 a_n11737_n15980.n11 a_n11737_n15980.n10 0.32719
R8846 a_n13990_8177.n62 a_n13990_8177.n60 7.94229
R8847 a_n13990_8177.n107 a_n13990_8177.n104 7.94229
R8848 a_n13990_8177.n253 a_n13990_8177.n251 7.22198
R8849 a_n13990_8177.n289 a_n13990_8177.n288 7.22198
R8850 a_n13990_8177.n238 a_n13990_8177.t144 6.77653
R8851 a_n13990_8177.n224 a_n13990_8177.t222 6.77653
R8852 a_n13990_8177.n230 a_n13990_8177.t272 6.7761
R8853 a_n13990_8177.n228 a_n13990_8177.t170 6.7761
R8854 a_n13990_8177.n21 a_n13990_8177.t182 6.77231
R8855 a_n13990_8177.n31 a_n13990_8177.t167 6.77231
R8856 a_n13990_8177.n215 a_n13990_8177.t292 6.58663
R8857 a_n13990_8177.n171 a_n13990_8177.t37 6.58663
R8858 a_n13990_8177.n355 a_n13990_8177.n354 6.50088
R8859 a_n13990_8177.n325 a_n13990_8177.n324 6.50088
R8860 a_n13990_8177.n216 a_n13990_8177.n213 5.95439
R8861 a_n13990_8177.n172 a_n13990_8177.n169 5.95439
R8862 a_n13990_8177.n59 a_n13990_8177.t213 5.69423
R8863 a_n13990_8177.n63 a_n13990_8177.t223 5.69423
R8864 a_n13990_8177.n106 a_n13990_8177.t108 5.69423
R8865 a_n13990_8177.n102 a_n13990_8177.t117 5.69423
R8866 a_n13990_8177.n242 a_n13990_8177.t237 5.50607
R8867 a_n13990_8177.n239 a_n13990_8177.t201 5.50607
R8868 a_n13990_8177.n269 a_n13990_8177.t135 5.50607
R8869 a_n13990_8177.n225 a_n13990_8177.t270 5.50607
R8870 a_n13990_8177.n241 a_n13990_8177.t121 5.50475
R8871 a_n13990_8177.n245 a_n13990_8177.t207 5.50475
R8872 a_n13990_8177.n246 a_n13990_8177.t150 5.50475
R8873 a_n13990_8177.n240 a_n13990_8177.t129 5.50475
R8874 a_n13990_8177.n268 a_n13990_8177.t197 5.50475
R8875 a_n13990_8177.n272 a_n13990_8177.t102 5.50475
R8876 a_n13990_8177.n273 a_n13990_8177.t228 5.50475
R8877 a_n13990_8177.n226 a_n13990_8177.t212 5.50475
R8878 a_n13990_8177.n59 a_n13990_8177.n58 5.49558
R8879 a_n13990_8177.n106 a_n13990_8177.n105 5.49558
R8880 a_n13990_8177.n213 a_n13990_8177.t53 5.31528
R8881 a_n13990_8177.n169 a_n13990_8177.t80 5.31528
R8882 a_n13990_8177.n359 a_n13990_8177.n357 4.92758
R8883 a_n13990_8177.n300 a_n13990_8177.n298 4.92758
R8884 a_n13990_8177.n38 a_n13990_8177.n338 4.92217
R8885 a_n13990_8177.n45 a_n13990_8177.n305 4.92217
R8886 a_n13990_8177.n0 a_n13990_8177.n99 4.22068
R8887 a_n13990_8177.t163 a_n13990_8177.n1 5.69068
R8888 a_n13990_8177.n98 a_n13990_8177.n2 4.22068
R8889 a_n13990_8177.n3 a_n13990_8177.n56 4.22068
R8890 a_n13990_8177.n4 a_n13990_8177.t149 5.69068
R8891 a_n13990_8177.n5 a_n13990_8177.n55 4.22068
R8892 a_n13990_8177.n7 a_n13990_8177.n132 3.84173
R8893 a_n13990_8177.n10 a_n13990_8177.n128 3.84173
R8894 a_n13990_8177.n346 a_n13990_8177.n32 3.65107
R8895 a_n13990_8177.n345 a_n13990_8177.n33 3.65107
R8896 a_n13990_8177.n344 a_n13990_8177.n34 3.65107
R8897 a_n13990_8177.n343 a_n13990_8177.n35 3.65107
R8898 a_n13990_8177.n341 a_n13990_8177.n36 3.65107
R8899 a_n13990_8177.n340 a_n13990_8177.n37 3.65107
R8900 a_n13990_8177.n339 a_n13990_8177.n38 3.65107
R8901 a_n13990_8177.n39 a_n13990_8177.n312 3.65107
R8902 a_n13990_8177.n40 a_n13990_8177.n311 3.65107
R8903 a_n13990_8177.n41 a_n13990_8177.n310 3.65107
R8904 a_n13990_8177.n42 a_n13990_8177.n309 3.65107
R8905 a_n13990_8177.n308 a_n13990_8177.n43 3.65107
R8906 a_n13990_8177.n307 a_n13990_8177.n44 3.65107
R8907 a_n13990_8177.n306 a_n13990_8177.n45 3.65107
R8908 a_n13990_8177.n12 a_n13990_8177.n380 4.0312
R8909 a_n13990_8177.t131 a_n13990_8177.n13 5.5012
R8910 a_n13990_8177.t206 a_n13990_8177.n14 5.5012
R8911 a_n13990_8177.n379 a_n13990_8177.n15 4.0312
R8912 a_n13990_8177.t164 a_n13990_8177.n16 5.5012
R8913 a_n13990_8177.t171 a_n13990_8177.n17 5.5012
R8914 a_n13990_8177.n378 a_n13990_8177.n18 4.0312
R8915 a_n13990_8177.t244 a_n13990_8177.n19 5.5012
R8916 a_n13990_8177.t269 a_n13990_8177.n20 5.5012
R8917 a_n13990_8177.n221 a_n13990_8177.n21 4.0312
R8918 a_n13990_8177.n22 a_n13990_8177.n263 4.0312
R8919 a_n13990_8177.t141 a_n13990_8177.n23 5.5012
R8920 a_n13990_8177.t263 a_n13990_8177.n24 5.5012
R8921 a_n13990_8177.n262 a_n13990_8177.n25 4.0312
R8922 a_n13990_8177.t226 a_n13990_8177.n26 5.5012
R8923 a_n13990_8177.t175 a_n13990_8177.n27 5.5012
R8924 a_n13990_8177.n261 a_n13990_8177.n28 4.0312
R8925 a_n13990_8177.t154 a_n13990_8177.n29 5.5012
R8926 a_n13990_8177.t224 a_n13990_8177.n30 5.5012
R8927 a_n13990_8177.n259 a_n13990_8177.n31 4.0312
R8928 a_n13990_8177.n6 a_n13990_8177.t28 5.31173
R8929 a_n13990_8177.n8 a_n13990_8177.t35 5.31173
R8930 a_n13990_8177.n9 a_n13990_8177.t26 5.31173
R8931 a_n13990_8177.n11 a_n13990_8177.t78 5.31173
R8932 a_n13990_8177.n212 a_n13990_8177.n210 4.50663
R8933 a_n13990_8177.n168 a_n13990_8177.n127 4.50663
R8934 a_n13990_8177.n133 a_n13990_8177.n8 4.46113
R8935 a_n13990_8177.n252 a_n13990_8177.t205 4.24002
R8936 a_n13990_8177.n232 a_n13990_8177.t217 4.24002
R8937 a_n13990_8177.n287 a_n13990_8177.t99 4.24002
R8938 a_n13990_8177.n278 a_n13990_8177.t214 4.24002
R8939 a_n13990_8177.n62 a_n13990_8177.n61 4.22423
R8940 a_n13990_8177.n104 a_n13990_8177.n103 4.22423
R8941 a_n13990_8177.n319 a_n13990_8177.t277 4.06712
R8942 a_n13990_8177.n317 a_n13990_8177.t52 4.06712
R8943 a_n13990_8177.n349 a_n13990_8177.t300 4.06712
R8944 a_n13990_8177.n295 a_n13990_8177.t72 4.06712
R8945 a_n13990_8177.n115 a_n13990_8177.t120 4.05054
R8946 a_n13990_8177.n120 a_n13990_8177.t147 4.05054
R8947 a_n13990_8177.n122 a_n13990_8177.t220 4.05054
R8948 a_n13990_8177.n109 a_n13990_8177.t180 4.05054
R8949 a_n13990_8177.n46 a_n13990_8177.t187 4.05054
R8950 a_n13990_8177.n392 a_n13990_8177.t264 4.05054
R8951 a_n13990_8177.n390 a_n13990_8177.t112 4.05054
R8952 a_n13990_8177.n48 a_n13990_8177.t199 4.05054
R8953 a_n13990_8177.n69 a_n13990_8177.t266 4.05054
R8954 a_n13990_8177.n74 a_n13990_8177.t116 4.05054
R8955 a_n13990_8177.n76 a_n13990_8177.t234 4.05054
R8956 a_n13990_8177.n83 a_n13990_8177.t202 4.05054
R8957 a_n13990_8177.n85 a_n13990_8177.t146 4.05054
R8958 a_n13990_8177.n91 a_n13990_8177.t126 4.05054
R8959 a_n13990_8177.n93 a_n13990_8177.t194 4.05054
R8960 a_n13990_8177.n64 a_n13990_8177.t138 4.05054
R8961 a_n13990_8177.n230 a_n13990_8177.n229 4.03475
R8962 a_n13990_8177.n244 a_n13990_8177.n243 4.03475
R8963 a_n13990_8177.n248 a_n13990_8177.n247 4.03475
R8964 a_n13990_8177.n238 a_n13990_8177.n237 4.03475
R8965 a_n13990_8177.n228 a_n13990_8177.n227 4.03475
R8966 a_n13990_8177.n271 a_n13990_8177.n270 4.03475
R8967 a_n13990_8177.n275 a_n13990_8177.n274 4.03475
R8968 a_n13990_8177.n224 a_n13990_8177.n223 4.03475
R8969 a_n13990_8177.n350 a_n13990_8177.n348 3.96014
R8970 a_n13990_8177.n320 a_n13990_8177.n297 3.96014
R8971 a_n13990_8177.n115 a_n13990_8177.t151 3.87765
R8972 a_n13990_8177.n120 a_n13990_8177.t179 3.87765
R8973 a_n13990_8177.n122 a_n13990_8177.t122 3.87765
R8974 a_n13990_8177.n109 a_n13990_8177.t259 3.87765
R8975 a_n13990_8177.n46 a_n13990_8177.t215 3.87765
R8976 a_n13990_8177.n392 a_n13990_8177.t192 3.87765
R8977 a_n13990_8177.n390 a_n13990_8177.t250 3.87765
R8978 a_n13990_8177.n48 a_n13990_8177.t209 3.87765
R8979 a_n13990_8177.n69 a_n13990_8177.t253 3.87765
R8980 a_n13990_8177.n74 a_n13990_8177.t110 3.87765
R8981 a_n13990_8177.n76 a_n13990_8177.t229 3.87765
R8982 a_n13990_8177.n83 a_n13990_8177.t190 3.87765
R8983 a_n13990_8177.n85 a_n13990_8177.t134 3.87765
R8984 a_n13990_8177.n91 a_n13990_8177.t119 3.87765
R8985 a_n13990_8177.n93 a_n13990_8177.t185 3.87765
R8986 a_n13990_8177.n64 a_n13990_8177.t127 3.87765
R8987 a_n13990_8177.n319 a_n13990_8177.t307 3.86107
R8988 a_n13990_8177.n317 a_n13990_8177.t68 3.86107
R8989 a_n13990_8177.n349 a_n13990_8177.t299 3.86107
R8990 a_n13990_8177.n295 a_n13990_8177.t70 3.86107
R8991 a_n13990_8177.n215 a_n13990_8177.n214 3.84528
R8992 a_n13990_8177.n212 a_n13990_8177.n211 3.84528
R8993 a_n13990_8177.n171 a_n13990_8177.n170 3.84528
R8994 a_n13990_8177.n168 a_n13990_8177.n167 3.84528
R8995 a_n13990_8177.n204 a_n13990_8177.n200 3.79678
R8996 a_n13990_8177.n187 a_n13990_8177.n183 3.79678
R8997 a_n13990_8177.n145 a_n13990_8177.n141 3.79678
R8998 a_n13990_8177.n160 a_n13990_8177.n156 3.79678
R8999 a_n13990_8177.n361 a_n13990_8177.n359 3.79678
R9000 a_n13990_8177.n369 a_n13990_8177.n367 3.79678
R9001 a_n13990_8177.n302 a_n13990_8177.n300 3.79678
R9002 a_n13990_8177.n334 a_n13990_8177.n332 3.79678
R9003 a_n13990_8177.n176 a_n13990_8177.n11 3.87644
R9004 a_n13990_8177.n196 a_n13990_8177.n192 3.73034
R9005 a_n13990_8177.n165 a_n13990_8177.n149 3.73034
R9006 a_n13990_8177.n252 a_n13990_8177.t193 3.68818
R9007 a_n13990_8177.n232 a_n13990_8177.t210 3.68818
R9008 a_n13990_8177.n287 a_n13990_8177.t265 3.68818
R9009 a_n13990_8177.n278 a_n13990_8177.t104 3.68818
R9010 a_n13990_8177.n365 a_n13990_8177.n364 3.65581
R9011 a_n13990_8177.n367 a_n13990_8177.n366 3.65581
R9012 a_n13990_8177.n369 a_n13990_8177.n368 3.65581
R9013 a_n13990_8177.n371 a_n13990_8177.n370 3.65581
R9014 a_n13990_8177.n363 a_n13990_8177.n362 3.65581
R9015 a_n13990_8177.n361 a_n13990_8177.n360 3.65581
R9016 a_n13990_8177.n359 a_n13990_8177.n358 3.65581
R9017 a_n13990_8177.n336 a_n13990_8177.n335 3.65581
R9018 a_n13990_8177.n334 a_n13990_8177.n333 3.65581
R9019 a_n13990_8177.n332 a_n13990_8177.n331 3.65581
R9020 a_n13990_8177.n330 a_n13990_8177.n329 3.65581
R9021 a_n13990_8177.n304 a_n13990_8177.n303 3.65581
R9022 a_n13990_8177.n302 a_n13990_8177.n301 3.65581
R9023 a_n13990_8177.n300 a_n13990_8177.n299 3.65581
R9024 a_n13990_8177.n372 a_n13990_8177.n371 3.64443
R9025 a_n13990_8177.n330 a_n13990_8177.n328 3.64443
R9026 a_n13990_8177.n35 a_n13990_8177.n342 3.64223
R9027 a_n13990_8177.n313 a_n13990_8177.n42 3.64223
R9028 a_n13990_8177.n96 a_n13990_8177.n63 3.25667
R9029 a_n13990_8177.n258 a_n13990_8177.n257 3.23904
R9030 a_n13990_8177.n286 a_n13990_8177.n220 3.23904
R9031 a_n13990_8177.n2 a_n13990_8177.n97 3.15553
R9032 a_n13990_8177.n387 a_n13990_8177.n5 3.15553
R9033 a_n13990_8177.n216 a_n13990_8177.n215 3.00663
R9034 a_n13990_8177.n172 a_n13990_8177.n171 3.00663
R9035 a_n13990_8177.n179 a_n13990_8177.n177 2.7866
R9036 a_n13990_8177.n182 a_n13990_8177.n180 2.7866
R9037 a_n13990_8177.n186 a_n13990_8177.n184 2.7866
R9038 a_n13990_8177.n190 a_n13990_8177.n188 2.7866
R9039 a_n13990_8177.n195 a_n13990_8177.n193 2.7866
R9040 a_n13990_8177.n199 a_n13990_8177.n197 2.7866
R9041 a_n13990_8177.n203 a_n13990_8177.n201 2.7866
R9042 a_n13990_8177.n207 a_n13990_8177.n205 2.7866
R9043 a_n13990_8177.n152 a_n13990_8177.n150 2.7866
R9044 a_n13990_8177.n155 a_n13990_8177.n153 2.7866
R9045 a_n13990_8177.n159 a_n13990_8177.n157 2.7866
R9046 a_n13990_8177.n163 a_n13990_8177.n161 2.7866
R9047 a_n13990_8177.n148 a_n13990_8177.n146 2.7866
R9048 a_n13990_8177.n144 a_n13990_8177.n142 2.7866
R9049 a_n13990_8177.n140 a_n13990_8177.n138 2.7866
R9050 a_n13990_8177.n136 a_n13990_8177.n134 2.7866
R9051 a_n13990_8177.n256 a_n13990_8177.n255 2.77002
R9052 a_n13990_8177.n235 a_n13990_8177.n234 2.77002
R9053 a_n13990_8177.n285 a_n13990_8177.n284 2.77002
R9054 a_n13990_8177.n281 a_n13990_8177.n280 2.77002
R9055 a_n13990_8177.n68 a_n13990_8177.n64 2.73714
R9056 a_n13990_8177.n236 a_n13990_8177.n232 2.73714
R9057 a_n13990_8177.n282 a_n13990_8177.n278 2.73714
R9058 a_n13990_8177.n296 a_n13990_8177.n294 2.73714
R9059 a_n13990_8177.n318 a_n13990_8177.n316 2.73714
R9060 a_n13990_8177.n52 a_n13990_8177.n48 2.73714
R9061 a_n13990_8177.n119 a_n13990_8177.n115 2.73672
R9062 a_n13990_8177.n73 a_n13990_8177.n69 2.73672
R9063 a_n13990_8177.n183 a_n13990_8177.n179 2.73672
R9064 a_n13990_8177.n156 a_n13990_8177.n152 2.73672
R9065 a_n13990_8177.n86 a_n13990_8177.n84 2.60203
R9066 a_n13990_8177.n246 a_n13990_8177.n245 2.60203
R9067 a_n13990_8177.n273 a_n13990_8177.n272 2.60203
R9068 a_n13990_8177.n110 a_n13990_8177.n47 2.60203
R9069 a_n13990_8177.n323 a_n13990_8177.n321 2.59712
R9070 a_n13990_8177.n316 a_n13990_8177.n314 2.59712
R9071 a_n13990_8177.n353 a_n13990_8177.n351 2.59712
R9072 a_n13990_8177.n294 a_n13990_8177.n292 2.59712
R9073 a_n13990_8177.n118 a_n13990_8177.n117 2.58054
R9074 a_n13990_8177.n113 a_n13990_8177.n112 2.58054
R9075 a_n13990_8177.n51 a_n13990_8177.n50 2.58054
R9076 a_n13990_8177.n72 a_n13990_8177.n71 2.58054
R9077 a_n13990_8177.n81 a_n13990_8177.n80 2.58054
R9078 a_n13990_8177.n89 a_n13990_8177.n88 2.58054
R9079 a_n13990_8177.n67 a_n13990_8177.n66 2.58054
R9080 a_n13990_8177.n397 a_n13990_8177.n396 2.58054
R9081 a_n13990_8177.n94 a_n13990_8177.n92 2.53418
R9082 a_n13990_8177.n77 a_n13990_8177.n75 2.53418
R9083 a_n13990_8177.n393 a_n13990_8177.n391 2.53418
R9084 a_n13990_8177.n123 a_n13990_8177.n121 2.53418
R9085 a_n13990_8177.n240 a_n13990_8177.n239 2.52436
R9086 a_n13990_8177.n242 a_n13990_8177.n241 2.52436
R9087 a_n13990_8177.n226 a_n13990_8177.n225 2.52436
R9088 a_n13990_8177.n269 a_n13990_8177.n268 2.52436
R9089 a_n13990_8177.n102 a_n13990_8177.n53 2.51873
R9090 a_n13990_8177.n355 a_n13990_8177.n296 2.46014
R9091 a_n13990_8177.n325 a_n13990_8177.n318 2.46014
R9092 a_n13990_8177.n118 a_n13990_8177.n116 2.40765
R9093 a_n13990_8177.n113 a_n13990_8177.n111 2.40765
R9094 a_n13990_8177.n51 a_n13990_8177.n49 2.40765
R9095 a_n13990_8177.n72 a_n13990_8177.n70 2.40765
R9096 a_n13990_8177.n81 a_n13990_8177.n79 2.40765
R9097 a_n13990_8177.n89 a_n13990_8177.n87 2.40765
R9098 a_n13990_8177.n67 a_n13990_8177.n65 2.40765
R9099 a_n13990_8177.n396 a_n13990_8177.n395 2.40765
R9100 a_n13990_8177.n323 a_n13990_8177.n322 2.39107
R9101 a_n13990_8177.n316 a_n13990_8177.n315 2.39107
R9102 a_n13990_8177.n353 a_n13990_8177.n352 2.39107
R9103 a_n13990_8177.n294 a_n13990_8177.n293 2.39107
R9104 a_n13990_8177.n175 a_n13990_8177.n9 2.37644
R9105 a_n13990_8177.n131 a_n13990_8177.n6 2.37644
R9106 a_n13990_8177.n60 a_n13990_8177.n57 2.23844
R9107 a_n13990_8177.n256 a_n13990_8177.n254 2.21818
R9108 a_n13990_8177.n235 a_n13990_8177.n233 2.21818
R9109 a_n13990_8177.n285 a_n13990_8177.n283 2.21818
R9110 a_n13990_8177.n281 a_n13990_8177.n279 2.21818
R9111 a_n13990_8177.n179 a_n13990_8177.n178 2.2016
R9112 a_n13990_8177.n182 a_n13990_8177.n181 2.2016
R9113 a_n13990_8177.n186 a_n13990_8177.n185 2.2016
R9114 a_n13990_8177.n190 a_n13990_8177.n189 2.2016
R9115 a_n13990_8177.n195 a_n13990_8177.n194 2.2016
R9116 a_n13990_8177.n199 a_n13990_8177.n198 2.2016
R9117 a_n13990_8177.n203 a_n13990_8177.n202 2.2016
R9118 a_n13990_8177.n207 a_n13990_8177.n206 2.2016
R9119 a_n13990_8177.n152 a_n13990_8177.n151 2.2016
R9120 a_n13990_8177.n155 a_n13990_8177.n154 2.2016
R9121 a_n13990_8177.n159 a_n13990_8177.n158 2.2016
R9122 a_n13990_8177.n163 a_n13990_8177.n162 2.2016
R9123 a_n13990_8177.n148 a_n13990_8177.n147 2.2016
R9124 a_n13990_8177.n144 a_n13990_8177.n143 2.2016
R9125 a_n13990_8177.n140 a_n13990_8177.n139 2.2016
R9126 a_n13990_8177.n136 a_n13990_8177.n135 2.2016
R9127 a_n13990_8177.n250 a_n13990_8177.n249 2.13841
R9128 a_n13990_8177.n258 a_n13990_8177.n231 2.13841
R9129 a_n13990_8177.n166 a_n13990_8177.n131 2.0852
R9130 a_n13990_8177.n326 a_n13990_8177.n313 2.0852
R9131 a_n13990_8177.n383 a_n13990_8177.n219 1.95191
R9132 a_n13990_8177.n210 a_n13990_8177.n54 1.90397
R9133 a_n13990_8177.n384 a_n13990_8177.n383 1.80854
R9134 a_n13990_8177.n375 a_n13990_8177.n54 1.80603
R9135 a_n13990_8177.n251 a_n13990_8177.n236 1.73904
R9136 a_n13990_8177.n289 a_n13990_8177.n282 1.73904
R9137 a_n13990_8177.n365 a_n13990_8177.n219 1.73609
R9138 a_n13990_8177.n337 a_n13990_8177.n336 1.73609
R9139 a_n13990_8177.n209 a_n13990_8177.n208 1.65018
R9140 a_n13990_8177.n137 a_n13990_8177.n133 1.65018
R9141 a_n13990_8177.n374 a_n13990_8177.n218 1.56167
R9142 a_n13990_8177.n100 a_n13990_8177.n0 1.65553
R9143 a_n13990_8177.n386 a_n13990_8177.n3 1.65553
R9144 a_n13990_8177.n96 a_n13990_8177.n95 1.5005
R9145 a_n13990_8177.n173 a_n13990_8177.n172 1.5005
R9146 a_n13990_8177.n175 a_n13990_8177.n174 1.5005
R9147 a_n13990_8177.n217 a_n13990_8177.n216 1.5005
R9148 a_n13990_8177.n166 a_n13990_8177.n165 1.5005
R9149 a_n13990_8177.n192 a_n13990_8177.n126 1.5005
R9150 a_n13990_8177.n290 a_n13990_8177.n289 1.5005
R9151 a_n13990_8177.n277 a_n13990_8177.n276 1.5005
R9152 a_n13990_8177.n260 a_n13990_8177.n222 1.5005
R9153 a_n13990_8177.n251 a_n13990_8177.n250 1.5005
R9154 a_n13990_8177.n377 a_n13990_8177.n376 1.5005
R9155 a_n13990_8177.n382 a_n13990_8177.n381 1.5005
R9156 a_n13990_8177.n267 a_n13990_8177.n266 1.5005
R9157 a_n13990_8177.n265 a_n13990_8177.n264 1.5005
R9158 a_n13990_8177.n356 a_n13990_8177.n355 1.5005
R9159 a_n13990_8177.n328 a_n13990_8177.n327 1.5005
R9160 a_n13990_8177.n342 a_n13990_8177.n291 1.5005
R9161 a_n13990_8177.n373 a_n13990_8177.n372 1.5005
R9162 a_n13990_8177.n326 a_n13990_8177.n325 1.5005
R9163 a_n13990_8177.n386 a_n13990_8177.n385 1.5005
R9164 a_n13990_8177.n108 a_n13990_8177.n107 1.5005
R9165 a_n13990_8177.n101 a_n13990_8177.n100 1.5005
R9166 a_n13990_8177.n78 a_n13990_8177.n57 1.5005
R9167 a_n13990_8177.n125 a_n13990_8177.n124 1.5005
R9168 a_n13990_8177.n389 a_n13990_8177.n388 1.5005
R9169 a_n13990_8177.n395 a_n13990_8177.t231 1.4705
R9170 a_n13990_8177.n395 a_n13990_8177.t172 1.4705
R9171 a_n13990_8177.n116 a_n13990_8177.t218 1.4705
R9172 a_n13990_8177.n116 a_n13990_8177.t159 1.4705
R9173 a_n13990_8177.n117 a_n13990_8177.t160 1.4705
R9174 a_n13990_8177.n117 a_n13990_8177.t235 1.4705
R9175 a_n13990_8177.n111 a_n13990_8177.t140 1.4705
R9176 a_n13990_8177.n111 a_n13990_8177.t236 1.4705
R9177 a_n13990_8177.n112 a_n13990_8177.t125 1.4705
R9178 a_n13990_8177.n112 a_n13990_8177.t268 1.4705
R9179 a_n13990_8177.n49 a_n13990_8177.t128 1.4705
R9180 a_n13990_8177.n49 a_n13990_8177.t247 1.4705
R9181 a_n13990_8177.n50 a_n13990_8177.t184 1.4705
R9182 a_n13990_8177.n50 a_n13990_8177.t174 1.4705
R9183 a_n13990_8177.n58 a_n13990_8177.t204 1.4705
R9184 a_n13990_8177.n58 a_n13990_8177.t258 1.4705
R9185 a_n13990_8177.n61 a_n13990_8177.t256 1.4705
R9186 a_n13990_8177.n61 a_n13990_8177.t137 1.4705
R9187 a_n13990_8177.n70 a_n13990_8177.t143 1.4705
R9188 a_n13990_8177.n70 a_n13990_8177.t262 1.4705
R9189 a_n13990_8177.n71 a_n13990_8177.t152 1.4705
R9190 a_n13990_8177.n71 a_n13990_8177.t98 1.4705
R9191 a_n13990_8177.n79 a_n13990_8177.t243 1.4705
R9192 a_n13990_8177.n79 a_n13990_8177.t169 1.4705
R9193 a_n13990_8177.n80 a_n13990_8177.t251 1.4705
R9194 a_n13990_8177.n80 a_n13990_8177.t178 1.4705
R9195 a_n13990_8177.n87 a_n13990_8177.t155 1.4705
R9196 a_n13990_8177.n87 a_n13990_8177.t101 1.4705
R9197 a_n13990_8177.n88 a_n13990_8177.t168 1.4705
R9198 a_n13990_8177.n88 a_n13990_8177.t113 1.4705
R9199 a_n13990_8177.n65 a_n13990_8177.t233 1.4705
R9200 a_n13990_8177.n65 a_n13990_8177.t181 1.4705
R9201 a_n13990_8177.n66 a_n13990_8177.t241 1.4705
R9202 a_n13990_8177.n66 a_n13990_8177.t191 1.4705
R9203 a_n13990_8177.n99 a_n13990_8177.t230 1.4705
R9204 a_n13990_8177.n99 a_n13990_8177.t225 1.4705
R9205 a_n13990_8177.n98 a_n13990_8177.t238 1.4705
R9206 a_n13990_8177.n98 a_n13990_8177.t107 1.4705
R9207 a_n13990_8177.n105 a_n13990_8177.t100 1.4705
R9208 a_n13990_8177.n105 a_n13990_8177.t156 1.4705
R9209 a_n13990_8177.n103 a_n13990_8177.t153 1.4705
R9210 a_n13990_8177.n103 a_n13990_8177.t216 1.4705
R9211 a_n13990_8177.n56 a_n13990_8177.t255 1.4705
R9212 a_n13990_8177.n56 a_n13990_8177.t132 1.4705
R9213 a_n13990_8177.n55 a_n13990_8177.t196 1.4705
R9214 a_n13990_8177.n55 a_n13990_8177.t208 1.4705
R9215 a_n13990_8177.n130 a_n13990_8177.t29 1.4705
R9216 a_n13990_8177.n130 a_n13990_8177.t321 1.4705
R9217 a_n13990_8177.n132 a_n13990_8177.t348 1.4705
R9218 a_n13990_8177.n132 a_n13990_8177.t342 1.4705
R9219 a_n13990_8177.n177 a_n13990_8177.t31 1.4705
R9220 a_n13990_8177.n177 a_n13990_8177.t288 1.4705
R9221 a_n13990_8177.n178 a_n13990_8177.t30 1.4705
R9222 a_n13990_8177.n178 a_n13990_8177.t351 1.4705
R9223 a_n13990_8177.n180 a_n13990_8177.t305 1.4705
R9224 a_n13990_8177.n180 a_n13990_8177.t79 1.4705
R9225 a_n13990_8177.n181 a_n13990_8177.t303 1.4705
R9226 a_n13990_8177.n181 a_n13990_8177.t336 1.4705
R9227 a_n13990_8177.n184 a_n13990_8177.t34 1.4705
R9228 a_n13990_8177.n184 a_n13990_8177.t7 1.4705
R9229 a_n13990_8177.n185 a_n13990_8177.t33 1.4705
R9230 a_n13990_8177.n185 a_n13990_8177.t15 1.4705
R9231 a_n13990_8177.n188 a_n13990_8177.t56 1.4705
R9232 a_n13990_8177.n188 a_n13990_8177.t349 1.4705
R9233 a_n13990_8177.n189 a_n13990_8177.t55 1.4705
R9234 a_n13990_8177.n189 a_n13990_8177.t320 1.4705
R9235 a_n13990_8177.n193 a_n13990_8177.t3 1.4705
R9236 a_n13990_8177.n193 a_n13990_8177.t344 1.4705
R9237 a_n13990_8177.n194 a_n13990_8177.t57 1.4705
R9238 a_n13990_8177.n194 a_n13990_8177.t86 1.4705
R9239 a_n13990_8177.n197 a_n13990_8177.t27 1.4705
R9240 a_n13990_8177.n197 a_n13990_8177.t32 1.4705
R9241 a_n13990_8177.n198 a_n13990_8177.t36 1.4705
R9242 a_n13990_8177.n198 a_n13990_8177.t40 1.4705
R9243 a_n13990_8177.n201 a_n13990_8177.t6 1.4705
R9244 a_n13990_8177.n201 a_n13990_8177.t44 1.4705
R9245 a_n13990_8177.n202 a_n13990_8177.t5 1.4705
R9246 a_n13990_8177.n202 a_n13990_8177.t43 1.4705
R9247 a_n13990_8177.n205 a_n13990_8177.t83 1.4705
R9248 a_n13990_8177.n205 a_n13990_8177.t54 1.4705
R9249 a_n13990_8177.n206 a_n13990_8177.t82 1.4705
R9250 a_n13990_8177.n206 a_n13990_8177.t346 1.4705
R9251 a_n13990_8177.n150 a_n13990_8177.t318 1.4705
R9252 a_n13990_8177.n150 a_n13990_8177.t347 1.4705
R9253 a_n13990_8177.n151 a_n13990_8177.t319 1.4705
R9254 a_n13990_8177.n151 a_n13990_8177.t350 1.4705
R9255 a_n13990_8177.n153 a_n13990_8177.t81 1.4705
R9256 a_n13990_8177.n153 a_n13990_8177.t84 1.4705
R9257 a_n13990_8177.n154 a_n13990_8177.t304 1.4705
R9258 a_n13990_8177.n154 a_n13990_8177.t85 1.4705
R9259 a_n13990_8177.n157 a_n13990_8177.t8 1.4705
R9260 a_n13990_8177.n157 a_n13990_8177.t39 1.4705
R9261 a_n13990_8177.n158 a_n13990_8177.t9 1.4705
R9262 a_n13990_8177.n158 a_n13990_8177.t41 1.4705
R9263 a_n13990_8177.n161 a_n13990_8177.t23 1.4705
R9264 a_n13990_8177.n161 a_n13990_8177.t289 1.4705
R9265 a_n13990_8177.n162 a_n13990_8177.t24 1.4705
R9266 a_n13990_8177.n162 a_n13990_8177.t290 1.4705
R9267 a_n13990_8177.n146 a_n13990_8177.t306 1.4705
R9268 a_n13990_8177.n146 a_n13990_8177.t343 1.4705
R9269 a_n13990_8177.n147 a_n13990_8177.t317 1.4705
R9270 a_n13990_8177.n147 a_n13990_8177.t345 1.4705
R9271 a_n13990_8177.n142 a_n13990_8177.t332 1.4705
R9272 a_n13990_8177.n142 a_n13990_8177.t10 1.4705
R9273 a_n13990_8177.n143 a_n13990_8177.t334 1.4705
R9274 a_n13990_8177.n143 a_n13990_8177.t11 1.4705
R9275 a_n13990_8177.n138 a_n13990_8177.t20 1.4705
R9276 a_n13990_8177.n138 a_n13990_8177.t17 1.4705
R9277 a_n13990_8177.n139 a_n13990_8177.t12 1.4705
R9278 a_n13990_8177.n139 a_n13990_8177.t18 1.4705
R9279 a_n13990_8177.n134 a_n13990_8177.t2 1.4705
R9280 a_n13990_8177.n134 a_n13990_8177.t45 1.4705
R9281 a_n13990_8177.n135 a_n13990_8177.t4 1.4705
R9282 a_n13990_8177.n135 a_n13990_8177.t46 1.4705
R9283 a_n13990_8177.n214 a_n13990_8177.t42 1.4705
R9284 a_n13990_8177.n214 a_n13990_8177.t333 1.4705
R9285 a_n13990_8177.n211 a_n13990_8177.t14 1.4705
R9286 a_n13990_8177.n211 a_n13990_8177.t25 1.4705
R9287 a_n13990_8177.n129 a_n13990_8177.t291 1.4705
R9288 a_n13990_8177.n129 a_n13990_8177.t21 1.4705
R9289 a_n13990_8177.n128 a_n13990_8177.t19 1.4705
R9290 a_n13990_8177.n128 a_n13990_8177.t335 1.4705
R9291 a_n13990_8177.n170 a_n13990_8177.t13 1.4705
R9292 a_n13990_8177.n170 a_n13990_8177.t16 1.4705
R9293 a_n13990_8177.n167 a_n13990_8177.t22 1.4705
R9294 a_n13990_8177.n167 a_n13990_8177.t38 1.4705
R9295 a_n13990_8177.n380 a_n13990_8177.t142 1.4705
R9296 a_n13990_8177.n380 a_n13990_8177.t227 1.4705
R9297 a_n13990_8177.n379 a_n13990_8177.t114 1.4705
R9298 a_n13990_8177.n379 a_n13990_8177.t248 1.4705
R9299 a_n13990_8177.n378 a_n13990_8177.t254 1.4705
R9300 a_n13990_8177.n378 a_n13990_8177.t162 1.4705
R9301 a_n13990_8177.n221 a_n13990_8177.t165 1.4705
R9302 a_n13990_8177.n221 a_n13990_8177.t157 1.4705
R9303 a_n13990_8177.n229 a_n13990_8177.t161 1.4705
R9304 a_n13990_8177.n229 a_n13990_8177.t105 1.4705
R9305 a_n13990_8177.n243 a_n13990_8177.t261 1.4705
R9306 a_n13990_8177.n243 a_n13990_8177.t186 1.4705
R9307 a_n13990_8177.n247 a_n13990_8177.t173 1.4705
R9308 a_n13990_8177.n247 a_n13990_8177.t115 1.4705
R9309 a_n13990_8177.n237 a_n13990_8177.t245 1.4705
R9310 a_n13990_8177.n237 a_n13990_8177.t198 1.4705
R9311 a_n13990_8177.n254 a_n13990_8177.t188 1.4705
R9312 a_n13990_8177.n254 a_n13990_8177.t240 1.4705
R9313 a_n13990_8177.n255 a_n13990_8177.t200 1.4705
R9314 a_n13990_8177.n255 a_n13990_8177.t249 1.4705
R9315 a_n13990_8177.n233 a_n13990_8177.t239 1.4705
R9316 a_n13990_8177.n233 a_n13990_8177.t124 1.4705
R9317 a_n13990_8177.n234 a_n13990_8177.t246 1.4705
R9318 a_n13990_8177.n234 a_n13990_8177.t130 1.4705
R9319 a_n13990_8177.n263 a_n13990_8177.t183 1.4705
R9320 a_n13990_8177.n263 a_n13990_8177.t123 1.4705
R9321 a_n13990_8177.n262 a_n13990_8177.t111 1.4705
R9322 a_n13990_8177.n262 a_n13990_8177.t211 1.4705
R9323 a_n13990_8177.n261 a_n13990_8177.t195 1.4705
R9324 a_n13990_8177.n261 a_n13990_8177.t133 1.4705
R9325 a_n13990_8177.n259 a_n13990_8177.t271 1.4705
R9326 a_n13990_8177.n259 a_n13990_8177.t219 1.4705
R9327 a_n13990_8177.n227 a_n13990_8177.t232 1.4705
R9328 a_n13990_8177.n227 a_n13990_8177.t176 1.4705
R9329 a_n13990_8177.n270 a_n13990_8177.t158 1.4705
R9330 a_n13990_8177.n270 a_n13990_8177.t252 1.4705
R9331 a_n13990_8177.n274 a_n13990_8177.t242 1.4705
R9332 a_n13990_8177.n274 a_n13990_8177.t189 1.4705
R9333 a_n13990_8177.n223 a_n13990_8177.t145 1.4705
R9334 a_n13990_8177.n223 a_n13990_8177.t267 1.4705
R9335 a_n13990_8177.n283 a_n13990_8177.t257 1.4705
R9336 a_n13990_8177.n283 a_n13990_8177.t139 1.4705
R9337 a_n13990_8177.n284 a_n13990_8177.t148 1.4705
R9338 a_n13990_8177.n284 a_n13990_8177.t103 1.4705
R9339 a_n13990_8177.n279 a_n13990_8177.t136 1.4705
R9340 a_n13990_8177.n279 a_n13990_8177.t203 1.4705
R9341 a_n13990_8177.n280 a_n13990_8177.t221 1.4705
R9342 a_n13990_8177.n280 a_n13990_8177.t166 1.4705
R9343 a_n13990_8177.n321 a_n13990_8177.t297 1.4705
R9344 a_n13990_8177.n321 a_n13990_8177.t285 1.4705
R9345 a_n13990_8177.n322 a_n13990_8177.t283 1.4705
R9346 a_n13990_8177.n322 a_n13990_8177.t287 1.4705
R9347 a_n13990_8177.n314 a_n13990_8177.t340 1.4705
R9348 a_n13990_8177.n314 a_n13990_8177.t278 1.4705
R9349 a_n13990_8177.n315 a_n13990_8177.t293 1.4705
R9350 a_n13990_8177.n315 a_n13990_8177.t309 1.4705
R9351 a_n13990_8177.n364 a_n13990_8177.t339 1.4705
R9352 a_n13990_8177.n364 a_n13990_8177.t282 1.4705
R9353 a_n13990_8177.n366 a_n13990_8177.t58 1.4705
R9354 a_n13990_8177.n366 a_n13990_8177.t51 1.4705
R9355 a_n13990_8177.n368 a_n13990_8177.t93 1.4705
R9356 a_n13990_8177.n368 a_n13990_8177.t286 1.4705
R9357 a_n13990_8177.n370 a_n13990_8177.t326 1.4705
R9358 a_n13990_8177.n370 a_n13990_8177.t279 1.4705
R9359 a_n13990_8177.n362 a_n13990_8177.t312 1.4705
R9360 a_n13990_8177.n362 a_n13990_8177.t323 1.4705
R9361 a_n13990_8177.n360 a_n13990_8177.t298 1.4705
R9362 a_n13990_8177.n360 a_n13990_8177.t311 1.4705
R9363 a_n13990_8177.n358 a_n13990_8177.t48 1.4705
R9364 a_n13990_8177.n358 a_n13990_8177.t330 1.4705
R9365 a_n13990_8177.n357 a_n13990_8177.t65 1.4705
R9366 a_n13990_8177.n357 a_n13990_8177.t325 1.4705
R9367 a_n13990_8177.n346 a_n13990_8177.t94 1.4705
R9368 a_n13990_8177.n346 a_n13990_8177.t59 1.4705
R9369 a_n13990_8177.n345 a_n13990_8177.t73 1.4705
R9370 a_n13990_8177.n345 a_n13990_8177.t331 1.4705
R9371 a_n13990_8177.n344 a_n13990_8177.t329 1.4705
R9372 a_n13990_8177.n344 a_n13990_8177.t284 1.4705
R9373 a_n13990_8177.n343 a_n13990_8177.t341 1.4705
R9374 a_n13990_8177.n343 a_n13990_8177.t316 1.4705
R9375 a_n13990_8177.n341 a_n13990_8177.t63 1.4705
R9376 a_n13990_8177.n341 a_n13990_8177.t97 1.4705
R9377 a_n13990_8177.n340 a_n13990_8177.t61 1.4705
R9378 a_n13990_8177.n340 a_n13990_8177.t75 1.4705
R9379 a_n13990_8177.n339 a_n13990_8177.t275 1.4705
R9380 a_n13990_8177.n339 a_n13990_8177.t315 1.4705
R9381 a_n13990_8177.n338 a_n13990_8177.t95 1.4705
R9382 a_n13990_8177.n338 a_n13990_8177.t76 1.4705
R9383 a_n13990_8177.n335 a_n13990_8177.t276 1.4705
R9384 a_n13990_8177.n335 a_n13990_8177.t308 1.4705
R9385 a_n13990_8177.n333 a_n13990_8177.t281 1.4705
R9386 a_n13990_8177.n333 a_n13990_8177.t50 1.4705
R9387 a_n13990_8177.n331 a_n13990_8177.t322 1.4705
R9388 a_n13990_8177.n331 a_n13990_8177.t338 1.4705
R9389 a_n13990_8177.n329 a_n13990_8177.t77 1.4705
R9390 a_n13990_8177.n329 a_n13990_8177.t96 1.4705
R9391 a_n13990_8177.n303 a_n13990_8177.t327 1.4705
R9392 a_n13990_8177.n303 a_n13990_8177.t69 1.4705
R9393 a_n13990_8177.n301 a_n13990_8177.t0 1.4705
R9394 a_n13990_8177.n301 a_n13990_8177.t314 1.4705
R9395 a_n13990_8177.n299 a_n13990_8177.t91 1.4705
R9396 a_n13990_8177.n299 a_n13990_8177.t90 1.4705
R9397 a_n13990_8177.n298 a_n13990_8177.t60 1.4705
R9398 a_n13990_8177.n298 a_n13990_8177.t337 1.4705
R9399 a_n13990_8177.n312 a_n13990_8177.t47 1.4705
R9400 a_n13990_8177.n312 a_n13990_8177.t280 1.4705
R9401 a_n13990_8177.n311 a_n13990_8177.t71 1.4705
R9402 a_n13990_8177.n311 a_n13990_8177.t67 1.4705
R9403 a_n13990_8177.n310 a_n13990_8177.t74 1.4705
R9404 a_n13990_8177.n310 a_n13990_8177.t310 1.4705
R9405 a_n13990_8177.n309 a_n13990_8177.t294 1.4705
R9406 a_n13990_8177.n309 a_n13990_8177.t328 1.4705
R9407 a_n13990_8177.n308 a_n13990_8177.t62 1.4705
R9408 a_n13990_8177.n308 a_n13990_8177.t324 1.4705
R9409 a_n13990_8177.n307 a_n13990_8177.t49 1.4705
R9410 a_n13990_8177.n307 a_n13990_8177.t88 1.4705
R9411 a_n13990_8177.n306 a_n13990_8177.t296 1.4705
R9412 a_n13990_8177.n306 a_n13990_8177.t295 1.4705
R9413 a_n13990_8177.n305 a_n13990_8177.t313 1.4705
R9414 a_n13990_8177.n305 a_n13990_8177.t274 1.4705
R9415 a_n13990_8177.n351 a_n13990_8177.t302 1.4705
R9416 a_n13990_8177.n351 a_n13990_8177.t92 1.4705
R9417 a_n13990_8177.n352 a_n13990_8177.t301 1.4705
R9418 a_n13990_8177.n352 a_n13990_8177.t1 1.4705
R9419 a_n13990_8177.n292 a_n13990_8177.t66 1.4705
R9420 a_n13990_8177.n292 a_n13990_8177.t89 1.4705
R9421 a_n13990_8177.n293 a_n13990_8177.t64 1.4705
R9422 a_n13990_8177.n293 a_n13990_8177.t87 1.4705
R9423 a_n13990_8177.t273 a_n13990_8177.n397 1.4705
R9424 a_n13990_8177.n397 a_n13990_8177.t177 1.4705
R9425 a_n13990_8177.n119 a_n13990_8177.n118 1.46537
R9426 a_n13990_8177.n121 a_n13990_8177.n120 1.46537
R9427 a_n13990_8177.n114 a_n13990_8177.n113 1.46537
R9428 a_n13990_8177.n110 a_n13990_8177.n109 1.46537
R9429 a_n13990_8177.n47 a_n13990_8177.n46 1.46537
R9430 a_n13990_8177.n396 a_n13990_8177.n394 1.46537
R9431 a_n13990_8177.n393 a_n13990_8177.n392 1.46537
R9432 a_n13990_8177.n52 a_n13990_8177.n51 1.46537
R9433 a_n13990_8177.n73 a_n13990_8177.n72 1.46537
R9434 a_n13990_8177.n75 a_n13990_8177.n74 1.46537
R9435 a_n13990_8177.n82 a_n13990_8177.n81 1.46537
R9436 a_n13990_8177.n84 a_n13990_8177.n83 1.46537
R9437 a_n13990_8177.n86 a_n13990_8177.n85 1.46537
R9438 a_n13990_8177.n90 a_n13990_8177.n89 1.46537
R9439 a_n13990_8177.n92 a_n13990_8177.n91 1.46537
R9440 a_n13990_8177.n68 a_n13990_8177.n67 1.46537
R9441 a_n13990_8177.n257 a_n13990_8177.n256 1.46537
R9442 a_n13990_8177.n253 a_n13990_8177.n252 1.46537
R9443 a_n13990_8177.n236 a_n13990_8177.n235 1.46537
R9444 a_n13990_8177.n286 a_n13990_8177.n285 1.46537
R9445 a_n13990_8177.n288 a_n13990_8177.n287 1.46537
R9446 a_n13990_8177.n282 a_n13990_8177.n281 1.46537
R9447 a_n13990_8177.n320 a_n13990_8177.n319 1.46537
R9448 a_n13990_8177.n324 a_n13990_8177.n323 1.46537
R9449 a_n13990_8177.n318 a_n13990_8177.n317 1.46537
R9450 a_n13990_8177.n350 a_n13990_8177.n349 1.46537
R9451 a_n13990_8177.n354 a_n13990_8177.n353 1.46537
R9452 a_n13990_8177.n296 a_n13990_8177.n295 1.46537
R9453 a_n13990_8177.n183 a_n13990_8177.n182 1.46537
R9454 a_n13990_8177.n187 a_n13990_8177.n186 1.46537
R9455 a_n13990_8177.n191 a_n13990_8177.n190 1.46537
R9456 a_n13990_8177.n196 a_n13990_8177.n195 1.46537
R9457 a_n13990_8177.n200 a_n13990_8177.n199 1.46537
R9458 a_n13990_8177.n204 a_n13990_8177.n203 1.46537
R9459 a_n13990_8177.n208 a_n13990_8177.n207 1.46537
R9460 a_n13990_8177.n156 a_n13990_8177.n155 1.46537
R9461 a_n13990_8177.n160 a_n13990_8177.n159 1.46537
R9462 a_n13990_8177.n164 a_n13990_8177.n163 1.46537
R9463 a_n13990_8177.n149 a_n13990_8177.n148 1.46537
R9464 a_n13990_8177.n145 a_n13990_8177.n144 1.46537
R9465 a_n13990_8177.n141 a_n13990_8177.n140 1.46537
R9466 a_n13990_8177.n137 a_n13990_8177.n136 1.46537
R9467 a_n13990_8177.n123 a_n13990_8177.n122 1.46535
R9468 a_n13990_8177.n391 a_n13990_8177.n390 1.46535
R9469 a_n13990_8177.n77 a_n13990_8177.n76 1.46535
R9470 a_n13990_8177.n94 a_n13990_8177.n93 1.46535
R9471 a_n13990_8177.n374 a_n13990_8177.n373 1.34705
R9472 a_n13990_8177.n218 a_n13990_8177.n217 1.2981
R9473 a_n13990_8177.n385 a_n13990_8177.n384 1.27763
R9474 a_n13990_8177.n394 a_n13990_8177.n47 1.27228
R9475 a_n13990_8177.n63 a_n13990_8177.n62 1.27228
R9476 a_n13990_8177.n92 a_n13990_8177.n90 1.27228
R9477 a_n13990_8177.n90 a_n13990_8177.n86 1.27228
R9478 a_n13990_8177.n84 a_n13990_8177.n82 1.27228
R9479 a_n13990_8177.n75 a_n13990_8177.n73 1.27228
R9480 a_n13990_8177.n104 a_n13990_8177.n102 1.27228
R9481 a_n13990_8177.n248 a_n13990_8177.n246 1.27228
R9482 a_n13990_8177.n245 a_n13990_8177.n244 1.27228
R9483 a_n13990_8177.n257 a_n13990_8177.n253 1.27228
R9484 a_n13990_8177.n275 a_n13990_8177.n273 1.27228
R9485 a_n13990_8177.n272 a_n13990_8177.n271 1.27228
R9486 a_n13990_8177.n288 a_n13990_8177.n286 1.27228
R9487 a_n13990_8177.n394 a_n13990_8177.n393 1.27228
R9488 a_n13990_8177.n114 a_n13990_8177.n110 1.27228
R9489 a_n13990_8177.n121 a_n13990_8177.n119 1.27228
R9490 a_n13990_8177.n208 a_n13990_8177.n204 1.27228
R9491 a_n13990_8177.n200 a_n13990_8177.n196 1.27228
R9492 a_n13990_8177.n191 a_n13990_8177.n187 1.27228
R9493 a_n13990_8177.n141 a_n13990_8177.n137 1.27228
R9494 a_n13990_8177.n149 a_n13990_8177.n145 1.27228
R9495 a_n13990_8177.n164 a_n13990_8177.n160 1.27228
R9496 a_n13990_8177.n213 a_n13990_8177.n212 1.27228
R9497 a_n13990_8177.n169 a_n13990_8177.n168 1.27228
R9498 a_n13990_8177.n363 a_n13990_8177.n361 1.27228
R9499 a_n13990_8177.n371 a_n13990_8177.n369 1.27228
R9500 a_n13990_8177.n367 a_n13990_8177.n365 1.27228
R9501 a_n13990_8177.n304 a_n13990_8177.n302 1.27228
R9502 a_n13990_8177.n332 a_n13990_8177.n330 1.27228
R9503 a_n13990_8177.n336 a_n13990_8177.n334 1.27228
R9504 a_n13990_8177.n354 a_n13990_8177.n350 1.27228
R9505 a_n13990_8177.n324 a_n13990_8177.n320 1.27228
R9506 a_n13990_8177.n239 a_n13990_8177.n238 1.26756
R9507 a_n13990_8177.n244 a_n13990_8177.n242 1.26756
R9508 a_n13990_8177.n225 a_n13990_8177.n224 1.26756
R9509 a_n13990_8177.n271 a_n13990_8177.n269 1.26756
R9510 a_n13990_8177.n383 a_n13990_8177.n382 1.23567
R9511 a_n13990_8177.n376 a_n13990_8177.n375 1.23455
R9512 a_n13990_8177.n387 a_n13990_8177.n54 1.18682
R9513 a_n13990_8177.n60 a_n13990_8177.n59 1.01873
R9514 a_n13990_8177.n107 a_n13990_8177.n106 1.01873
R9515 a_n13990_8177.n327 a_n13990_8177.n291 0.822966
R9516 a_n13990_8177.n347 a_n13990_8177.n337 0.822966
R9517 a_n13990_8177.n249 a_n13990_8177.n240 0.796291
R9518 a_n13990_8177.n241 a_n13990_8177.n231 0.796291
R9519 a_n13990_8177.n276 a_n13990_8177.n226 0.796291
R9520 a_n13990_8177.n268 a_n13990_8177.n267 0.796291
R9521 a_n13990_8177.n250 a_n13990_8177.n222 0.780703
R9522 a_n13990_8177.n376 a_n13990_8177.n290 0.780703
R9523 a_n13990_8177.n265 a_n13990_8177.n258 0.780703
R9524 a_n13990_8177.n382 a_n13990_8177.n220 0.780703
R9525 a_n13990_8177.n97 a_n13990_8177.n96 0.778574
R9526 a_n13990_8177.n388 a_n13990_8177.n387 0.778574
R9527 a_n13990_8177.n101 a_n13990_8177.n57 0.778574
R9528 a_n13990_8177.n385 a_n13990_8177.n125 0.778574
R9529 a_n13990_8177.n388 a_n13990_8177.n53 0.738439
R9530 a_n13990_8177.n125 a_n13990_8177.n108 0.738439
R9531 a_n13990_8177.n210 a_n13990_8177.n209 0.737223
R9532 a_n13990_8177.n133 a_n13990_8177.n127 0.737223
R9533 a_n13990_8177.n217 a_n13990_8177.n126 0.737223
R9534 a_n13990_8177.n173 a_n13990_8177.n166 0.737223
R9535 a_n13990_8177.n176 a_n13990_8177.n127 0.725061
R9536 a_n13990_8177.n174 a_n13990_8177.n173 0.725061
R9537 a_n13990_8177.n95 a_n13990_8177.n94 0.699581
R9538 a_n13990_8177.n78 a_n13990_8177.n77 0.699581
R9539 a_n13990_8177.n391 a_n13990_8177.n389 0.699581
R9540 a_n13990_8177.n124 a_n13990_8177.n123 0.699581
R9541 a_n13990_8177.n373 a_n13990_8177.n356 0.639318
R9542 a_n13990_8177.n327 a_n13990_8177.n326 0.639318
R9543 a_n13990_8177.n348 a_n13990_8177.n219 0.639318
R9544 a_n13990_8177.n337 a_n13990_8177.n297 0.639318
R9545 a_n13990_8177.n290 a_n13990_8177.n277 0.638405
R9546 a_n13990_8177.n266 a_n13990_8177.n220 0.638405
R9547 a_n13990_8177.n277 a_n13990_8177.n222 0.628372
R9548 a_n13990_8177.n266 a_n13990_8177.n265 0.628372
R9549 a_n13990_8177.n375 a_n13990_8177.n374 0.606869
R9550 a_n13990_8177.n384 a_n13990_8177.n218 0.60536
R9551 a_n13990_8177.n209 a_n13990_8177.n176 0.585196
R9552 a_n13990_8177.n174 a_n13990_8177.n126 0.585196
R9553 a_n13990_8177.n356 a_n13990_8177.n291 0.585196
R9554 a_n13990_8177.n348 a_n13990_8177.n347 0.585196
R9555 a_n13990_8177.n95 a_n13990_8177.n68 0.557791
R9556 a_n13990_8177.n82 a_n13990_8177.n78 0.557791
R9557 a_n13990_8177.n389 a_n13990_8177.n52 0.557791
R9558 a_n13990_8177.n124 a_n13990_8177.n114 0.557791
R9559 a_n13990_8177.n97 a_n13990_8177.n53 0.530466
R9560 a_n13990_8177.n108 a_n13990_8177.n101 0.530466
R9561 a_n13990_8177.n249 a_n13990_8177.n248 0.476484
R9562 a_n13990_8177.n231 a_n13990_8177.n230 0.476484
R9563 a_n13990_8177.n276 a_n13990_8177.n275 0.476484
R9564 a_n13990_8177.n267 a_n13990_8177.n228 0.476484
R9565 a_n13990_8177.n28 a_n13990_8177.n260 0.478684
R9566 a_n13990_8177.n264 a_n13990_8177.n22 0.478684
R9567 a_n13990_8177.n18 a_n13990_8177.n377 0.478684
R9568 a_n13990_8177.n381 a_n13990_8177.n12 0.478684
R9569 a_n13990_8177.n372 a_n13990_8177.n363 0.236091
R9570 a_n13990_8177.n328 a_n13990_8177.n304 0.236091
R9571 a_n13990_8177.n192 a_n13990_8177.n191 0.150184
R9572 a_n13990_8177.n165 a_n13990_8177.n164 0.150184
R9573 a_n13990_8177.n1 a_n13990_8177.n2 1.27228
R9574 a_n13990_8177.n100 a_n13990_8177.n1 7.30549
R9575 a_n13990_8177.t109 a_n13990_8177.n0 6.96214
R9576 a_n13990_8177.n4 a_n13990_8177.n5 1.27228
R9577 a_n13990_8177.n386 a_n13990_8177.n4 7.30549
R9578 a_n13990_8177.t260 a_n13990_8177.n3 6.96214
R9579 a_n13990_8177.n10 a_n13990_8177.n11 1.26457
R9580 a_n13990_8177.n175 a_n13990_8177.n10 6.59229
R9581 a_n13990_8177.n129 a_n13990_8177.n9 5.10549
R9582 a_n13990_8177.n7 a_n13990_8177.n8 1.26457
R9583 a_n13990_8177.n131 a_n13990_8177.n7 6.59229
R9584 a_n13990_8177.n130 a_n13990_8177.n6 5.10549
R9585 a_n13990_8177.n30 a_n13990_8177.n31 1.27228
R9586 a_n13990_8177.n29 a_n13990_8177.n30 2.51878
R9587 a_n13990_8177.n260 a_n13990_8177.n29 0.794091
R9588 a_n13990_8177.n27 a_n13990_8177.n28 1.27228
R9589 a_n13990_8177.n26 a_n13990_8177.n27 2.60203
R9590 a_n13990_8177.n25 a_n13990_8177.n26 1.27228
R9591 a_n13990_8177.n24 a_n13990_8177.n25 1.27228
R9592 a_n13990_8177.n23 a_n13990_8177.n24 2.51878
R9593 a_n13990_8177.n264 a_n13990_8177.n23 0.794091
R9594 a_n13990_8177.t118 a_n13990_8177.n22 6.77266
R9595 a_n13990_8177.n20 a_n13990_8177.n21 1.27228
R9596 a_n13990_8177.n19 a_n13990_8177.n20 2.51878
R9597 a_n13990_8177.n377 a_n13990_8177.n19 0.794091
R9598 a_n13990_8177.n17 a_n13990_8177.n18 1.27228
R9599 a_n13990_8177.n16 a_n13990_8177.n17 2.60203
R9600 a_n13990_8177.n15 a_n13990_8177.n16 1.27228
R9601 a_n13990_8177.n14 a_n13990_8177.n15 1.27228
R9602 a_n13990_8177.n13 a_n13990_8177.n14 2.51878
R9603 a_n13990_8177.n381 a_n13990_8177.n13 0.794091
R9604 a_n13990_8177.t106 a_n13990_8177.n12 6.77266
R9605 a_n13990_8177.n37 a_n13990_8177.n38 3.79678
R9606 a_n13990_8177.n36 a_n13990_8177.n37 1.27228
R9607 a_n13990_8177.n342 a_n13990_8177.n36 0.238291
R9608 a_n13990_8177.n34 a_n13990_8177.n35 1.27228
R9609 a_n13990_8177.n33 a_n13990_8177.n34 3.79678
R9610 a_n13990_8177.n32 a_n13990_8177.n33 1.27228
R9611 a_n13990_8177.n347 a_n13990_8177.n32 1.73829
R9612 a_n13990_8177.n44 a_n13990_8177.n45 3.79678
R9613 a_n13990_8177.n43 a_n13990_8177.n44 1.27228
R9614 a_n13990_8177.n313 a_n13990_8177.n43 0.238291
R9615 a_n13990_8177.n41 a_n13990_8177.n42 1.27228
R9616 a_n13990_8177.n40 a_n13990_8177.n41 3.79678
R9617 a_n13990_8177.n39 a_n13990_8177.n40 1.27228
R9618 a_n13990_8177.n297 a_n13990_8177.n39 2.32299
R9619 a_n11317_n20927.t1 a_n11317_n20927.t5 23.2164
R9620 a_n11317_n20927.t4 a_n11317_n20927.t1 17.4491
R9621 a_n11317_n20927.t1 a_n11317_n20927.t3 17.1874
R9622 a_n11317_n20927.t0 a_n11317_n20927.t1 16.5634
R9623 VP.n11 VP.t25 8.38704
R9624 VP.n311 VP.t69 8.38704
R9625 VP.n125 VP.t7 8.37857
R9626 VP.n248 VP.t19 8.37857
R9627 VP.n58 VP.t60 8.31301
R9628 VP.n209 VP.t85 8.31301
R9629 VP.n388 VP.t5 8.29322
R9630 VP.n147 VP.t84 8.29322
R9631 VP.n387 VP.t3 8.10567
R9632 VP.n385 VP.t62 8.10567
R9633 VP.n384 VP.t81 8.10567
R9634 VP.n0 VP.t18 8.10567
R9635 VP.n339 VP.t47 8.10567
R9636 VP.n340 VP.t43 8.10567
R9637 VP.n322 VP.t40 8.10567
R9638 VP.n316 VP.t41 8.10567
R9639 VP.n310 VP.t13 8.10567
R9640 VP.n326 VP.t78 8.10567
R9641 VP.n325 VP.t20 8.10567
R9642 VP.n324 VP.t38 8.10567
R9643 VP.n332 VP.t65 8.10567
R9644 VP.n331 VP.t87 8.10567
R9645 VP.n369 VP.t54 8.10567
R9646 VP.n375 VP.t74 8.10567
R9647 VP.n116 VP.t46 8.10567
R9648 VP.n109 VP.t23 8.10567
R9649 VP.n103 VP.t4 8.10567
R9650 VP.n97 VP.t67 8.10567
R9651 VP.n120 VP.t30 8.10567
R9652 VP.n119 VP.t2 8.10567
R9653 VP.n118 VP.t32 8.10567
R9654 VP.n124 VP.t35 8.10567
R9655 VP.n123 VP.t76 8.10567
R9656 VP.n135 VP.t83 8.10567
R9657 VP.n53 VP.t11 8.10567
R9658 VP.n62 VP.t73 8.10567
R9659 VP.n57 VP.t66 8.10567
R9660 VP.n75 VP.t82 8.10567
R9661 VP.n74 VP.t55 8.10567
R9662 VP.n73 VP.t61 8.10567
R9663 VP.n95 VP.t64 8.10567
R9664 VP.n88 VP.t68 8.10567
R9665 VP.n81 VP.t22 8.10567
R9666 VP.n52 VP.t28 8.10567
R9667 VP.n39 VP.t44 8.10567
R9668 VP.n37 VP.t10 8.10567
R9669 VP.n36 VP.t72 8.10567
R9670 VP.n180 VP.t37 8.10567
R9671 VP.n161 VP.t29 8.10567
R9672 VP.n162 VP.t0 8.10567
R9673 VP.n163 VP.t31 8.10567
R9674 VP.n146 VP.t24 8.10567
R9675 VP.n144 VP.t12 8.10567
R9676 VP.n143 VP.t48 8.10567
R9677 VP.n22 VP.t71 8.10567
R9678 VP.n16 VP.t14 8.10567
R9679 VP.n10 VP.t51 8.10567
R9680 VP.n26 VP.t80 8.10567
R9681 VP.n25 VP.t53 8.10567
R9682 VP.n24 VP.t59 8.10567
R9683 VP.n32 VP.t27 8.10567
R9684 VP.n31 VP.t58 8.10567
R9685 VP.n192 VP.t50 8.10567
R9686 VP.n198 VP.t86 8.10567
R9687 VP.n242 VP.t34 8.10567
R9688 VP.n238 VP.t63 8.10567
R9689 VP.n237 VP.t26 8.10567
R9690 VP.n281 VP.t52 8.10567
R9691 VP.n261 VP.t16 8.10567
R9692 VP.n262 VP.t45 8.10567
R9693 VP.n263 VP.t42 8.10567
R9694 VP.n247 VP.t15 8.10567
R9695 VP.n245 VP.t75 8.10567
R9696 VP.n243 VP.t6 8.10567
R9697 VP.n223 VP.t56 8.10567
R9698 VP.n216 VP.t57 8.10567
R9699 VP.n210 VP.t33 8.10567
R9700 VP.n227 VP.t77 8.10567
R9701 VP.n226 VP.t17 8.10567
R9702 VP.n225 VP.t36 8.10567
R9703 VP.n283 VP.t79 8.10567
R9704 VP.n231 VP.t8 8.10567
R9705 VP.n230 VP.t70 8.10567
R9706 VP.n300 VP.t1 8.10567
R9707 VP.n342 VP.t21 8.10567
R9708 VP.n337 VP.t49 8.10567
R9709 VP.n336 VP.t9 8.10567
R9710 VP.n357 VP.t39 8.10567
R9711 VP.n381 VP.n380 7.37198
R9712 VP.n359 VP.n332 4.64261
R9713 VP.n182 VP.n32 4.64261
R9714 VP.n96 VP.n95 4.61892
R9715 VP.n284 VP.n283 4.61892
R9716 VP.n98 VP.n97 4.61655
R9717 VP.n282 VP.n281 4.61655
R9718 VP.n60 VP.n59 4.5005
R9719 VP.n61 VP.n56 4.5005
R9720 VP.n64 VP.n63 4.5005
R9721 VP.n65 VP.n55 4.5005
R9722 VP.n67 VP.n66 4.5005
R9723 VP.n68 VP.n54 4.5005
R9724 VP.n70 VP.n69 4.5005
R9725 VP.n72 VP.n71 4.5005
R9726 VP.n77 VP.n76 4.5005
R9727 VP.n79 VP.n78 4.5005
R9728 VP.n80 VP.n51 4.5005
R9729 VP.n83 VP.n82 4.5005
R9730 VP.n84 VP.n50 4.5005
R9731 VP.n86 VP.n85 4.5005
R9732 VP.n87 VP.n49 4.5005
R9733 VP.n90 VP.n89 4.5005
R9734 VP.n91 VP.n48 4.5005
R9735 VP.n93 VP.n92 4.5005
R9736 VP.n94 VP.n47 4.5005
R9737 VP.n99 VP.n46 4.5005
R9738 VP.n101 VP.n100 4.5005
R9739 VP.n102 VP.n45 4.5005
R9740 VP.n105 VP.n104 4.5005
R9741 VP.n106 VP.n44 4.5005
R9742 VP.n108 VP.n107 4.5005
R9743 VP.n110 VP.n43 4.5005
R9744 VP.n112 VP.n111 4.5005
R9745 VP.n113 VP.n42 4.5005
R9746 VP.n115 VP.n114 4.5005
R9747 VP.n117 VP.n40 4.5005
R9748 VP.n137 VP.n136 4.5005
R9749 VP.n134 VP.n41 4.5005
R9750 VP.n133 VP.n132 4.5005
R9751 VP.n131 VP.n121 4.5005
R9752 VP.n130 VP.n129 4.5005
R9753 VP.n128 VP.n122 4.5005
R9754 VP.n127 VP.n126 4.5005
R9755 VP.n23 VP.n5 4.5005
R9756 VP.n21 VP.n20 4.5005
R9757 VP.n19 VP.n7 4.5005
R9758 VP.n18 VP.n17 4.5005
R9759 VP.n15 VP.n8 4.5005
R9760 VP.n14 VP.n13 4.5005
R9761 VP.n12 VP.n9 4.5005
R9762 VP.n201 VP.n200 4.5005
R9763 VP.n199 VP.n6 4.5005
R9764 VP.n197 VP.n196 4.5005
R9765 VP.n195 VP.n27 4.5005
R9766 VP.n194 VP.n193 4.5005
R9767 VP.n191 VP.n28 4.5005
R9768 VP.n190 VP.n189 4.5005
R9769 VP.n188 VP.n29 4.5005
R9770 VP.n187 VP.n186 4.5005
R9771 VP.n185 VP.n30 4.5005
R9772 VP.n184 VP.n183 4.5005
R9773 VP.n165 VP.n164 4.5005
R9774 VP.n167 VP.n166 4.5005
R9775 VP.n168 VP.n38 4.5005
R9776 VP.n170 VP.n169 4.5005
R9777 VP.n172 VP.n171 4.5005
R9778 VP.n173 VP.n35 4.5005
R9779 VP.n175 VP.n174 4.5005
R9780 VP.n176 VP.n34 4.5005
R9781 VP.n178 VP.n177 4.5005
R9782 VP.n179 VP.n33 4.5005
R9783 VP.n160 VP.n159 4.5005
R9784 VP.n158 VP.n141 4.5005
R9785 VP.n157 VP.n156 4.5005
R9786 VP.n155 VP.n142 4.5005
R9787 VP.n154 VP.n153 4.5005
R9788 VP.n152 VP.n151 4.5005
R9789 VP.n150 VP.n145 4.5005
R9790 VP.n149 VP.n148 4.5005
R9791 VP.n212 VP.n211 4.5005
R9792 VP.n213 VP.n208 4.5005
R9793 VP.n215 VP.n214 4.5005
R9794 VP.n217 VP.n207 4.5005
R9795 VP.n219 VP.n218 4.5005
R9796 VP.n220 VP.n206 4.5005
R9797 VP.n222 VP.n221 4.5005
R9798 VP.n224 VP.n204 4.5005
R9799 VP.n302 VP.n301 4.5005
R9800 VP.n299 VP.n205 4.5005
R9801 VP.n298 VP.n297 4.5005
R9802 VP.n296 VP.n228 4.5005
R9803 VP.n295 VP.n294 4.5005
R9804 VP.n293 VP.n229 4.5005
R9805 VP.n292 VP.n291 4.5005
R9806 VP.n290 VP.n289 4.5005
R9807 VP.n288 VP.n232 4.5005
R9808 VP.n287 VP.n286 4.5005
R9809 VP.n285 VP.n233 4.5005
R9810 VP.n280 VP.n234 4.5005
R9811 VP.n279 VP.n278 4.5005
R9812 VP.n277 VP.n235 4.5005
R9813 VP.n276 VP.n275 4.5005
R9814 VP.n274 VP.n236 4.5005
R9815 VP.n273 VP.n272 4.5005
R9816 VP.n271 VP.n270 4.5005
R9817 VP.n269 VP.n239 4.5005
R9818 VP.n268 VP.n267 4.5005
R9819 VP.n266 VP.n240 4.5005
R9820 VP.n265 VP.n264 4.5005
R9821 VP.n260 VP.n259 4.5005
R9822 VP.n258 VP.n257 4.5005
R9823 VP.n256 VP.n244 4.5005
R9824 VP.n255 VP.n254 4.5005
R9825 VP.n253 VP.n252 4.5005
R9826 VP.n251 VP.n246 4.5005
R9827 VP.n250 VP.n249 4.5005
R9828 VP.n323 VP.n305 4.5005
R9829 VP.n321 VP.n320 4.5005
R9830 VP.n319 VP.n307 4.5005
R9831 VP.n318 VP.n317 4.5005
R9832 VP.n315 VP.n308 4.5005
R9833 VP.n314 VP.n313 4.5005
R9834 VP.n312 VP.n309 4.5005
R9835 VP.n378 VP.n377 4.5005
R9836 VP.n376 VP.n306 4.5005
R9837 VP.n374 VP.n373 4.5005
R9838 VP.n372 VP.n327 4.5005
R9839 VP.n371 VP.n370 4.5005
R9840 VP.n368 VP.n328 4.5005
R9841 VP.n367 VP.n366 4.5005
R9842 VP.n365 VP.n329 4.5005
R9843 VP.n364 VP.n363 4.5005
R9844 VP.n362 VP.n330 4.5005
R9845 VP.n361 VP.n360 4.5005
R9846 VP.n341 VP.n2 4.5005
R9847 VP.n344 VP.n343 4.5005
R9848 VP.n345 VP.n338 4.5005
R9849 VP.n347 VP.n346 4.5005
R9850 VP.n349 VP.n348 4.5005
R9851 VP.n350 VP.n335 4.5005
R9852 VP.n352 VP.n351 4.5005
R9853 VP.n353 VP.n334 4.5005
R9854 VP.n355 VP.n354 4.5005
R9855 VP.n356 VP.n333 4.5005
R9856 VP.n401 VP.n400 4.5005
R9857 VP.n399 VP.n1 4.5005
R9858 VP.n398 VP.n397 4.5005
R9859 VP.n396 VP.n383 4.5005
R9860 VP.n395 VP.n394 4.5005
R9861 VP.n393 VP.n392 4.5005
R9862 VP.n391 VP.n386 4.5005
R9863 VP.n390 VP.n389 4.5005
R9864 VP.n182 VP.n181 3.03856
R9865 VP.n359 VP.n358 3.03856
R9866 VP.n98 VP.n96 3.0245
R9867 VP.n284 VP.n282 3.0245
R9868 VP.n203 VP.n4 2.30989
R9869 VP.n139 VP.n138 2.30989
R9870 VP.n181 VP.n180 2.25752
R9871 VP.n358 VP.n357 2.25752
R9872 VP.n71 VP.n4 2.18975
R9873 VP.n138 VP.n40 2.18975
R9874 VP.n303 VP.n204 2.18975
R9875 VP.n265 VP.n241 2.18975
R9876 VP.n202 VP.n5 2.16725
R9877 VP.n165 VP.n140 2.16725
R9878 VP.n379 VP.n305 2.16725
R9879 VP.n382 VP.n2 2.16725
R9880 VP.n304 VP.n303 1.5005
R9881 VP.n203 VP.n202 1.5005
R9882 VP.n241 VP.n3 1.5005
R9883 VP.n140 VP.n139 1.5005
R9884 VP.n382 VP.n381 1.5005
R9885 VP.n380 VP.n379 1.5005
R9886 VP.n148 VP.n147 1.392
R9887 VP.n389 VP.n388 1.392
R9888 VP.n59 VP.n58 1.38741
R9889 VP.n212 VP.n209 1.38741
R9890 VP.n136 VP.n120 1.24866
R9891 VP.n76 VP.n75 1.24866
R9892 VP.n261 VP.n260 1.24866
R9893 VP.n301 VP.n227 1.24866
R9894 VP.n118 VP.n117 1.24629
R9895 VP.n73 VP.n72 1.24629
R9896 VP.n264 VP.n263 1.24629
R9897 VP.n225 VP.n224 1.24629
R9898 VP.n304 VP.n203 1.23709
R9899 VP.n139 VP.n3 1.23709
R9900 VP.n324 VP.n323 1.22261
R9901 VP.n164 VP.n163 1.22261
R9902 VP.n24 VP.n23 1.22261
R9903 VP.n341 VP.n340 1.22261
R9904 VP.n377 VP.n326 1.21313
R9905 VP.n161 VP.n160 1.21313
R9906 VP.n200 VP.n26 1.21313
R9907 VP.n12 VP.n11 1.12904
R9908 VP.n312 VP.n311 1.12904
R9909 VP.n126 VP.n125 1.11862
R9910 VP.n249 VP.n248 1.11862
R9911 VP VP.n0 1.06037
R9912 VP.n380 VP.n304 0.809892
R9913 VP.n381 VP.n3 0.809892
R9914 VP.n77 VP.n4 0.752
R9915 VP.n138 VP.n137 0.752
R9916 VP.n303 VP.n302 0.752
R9917 VP.n259 VP.n241 0.752
R9918 VP.n202 VP.n201 0.71825
R9919 VP.n159 VP.n140 0.71825
R9920 VP.n379 VP.n378 0.71825
R9921 VP.n400 VP.n382 0.71825
R9922 VP.n325 VP.n324 0.673132
R9923 VP.n326 VP.n325 0.673132
R9924 VP.n119 VP.n118 0.673132
R9925 VP.n120 VP.n119 0.673132
R9926 VP.n74 VP.n73 0.673132
R9927 VP.n75 VP.n74 0.673132
R9928 VP.n163 VP.n162 0.673132
R9929 VP.n162 VP.n161 0.673132
R9930 VP.n25 VP.n24 0.673132
R9931 VP.n26 VP.n25 0.673132
R9932 VP.n263 VP.n262 0.673132
R9933 VP.n262 VP.n261 0.673132
R9934 VP.n226 VP.n225 0.673132
R9935 VP.n227 VP.n226 0.673132
R9936 VP.n340 VP.n339 0.673132
R9937 VP.n339 VP.n0 0.673132
R9938 VP.n147 VP.n146 0.45279
R9939 VP.n388 VP.n387 0.45279
R9940 VP.n58 VP.n57 0.430924
R9941 VP.n210 VP.n209 0.430924
R9942 VP.n128 VP.n127 0.394842
R9943 VP.n108 VP.n44 0.394842
R9944 VP.n87 VP.n86 0.394842
R9945 VP.n63 VP.n61 0.394842
R9946 VP.n251 VP.n250 0.394842
R9947 VP.n274 VP.n273 0.394842
R9948 VP.n293 VP.n292 0.394842
R9949 VP.n215 VP.n208 0.394842
R9950 VP.n133 VP.n121 0.381816
R9951 VP.n102 VP.n101 0.381816
R9952 VP.n82 VP.n80 0.381816
R9953 VP.n256 VP.n255 0.381816
R9954 VP.n279 VP.n235 0.381816
R9955 VP.n298 VP.n228 0.381816
R9956 VP.n374 VP.n327 0.379447
R9957 VP.n368 VP.n367 0.379447
R9958 VP.n363 VP.n362 0.379447
R9959 VP.n314 VP.n309 0.379447
R9960 VP.n317 VP.n307 0.379447
R9961 VP.n156 VP.n155 0.379447
R9962 VP.n151 VP.n150 0.379447
R9963 VP.n179 VP.n178 0.379447
R9964 VP.n174 VP.n173 0.379447
R9965 VP.n169 VP.n168 0.379447
R9966 VP.n197 VP.n27 0.379447
R9967 VP.n191 VP.n190 0.379447
R9968 VP.n186 VP.n185 0.379447
R9969 VP.n14 VP.n9 0.379447
R9970 VP.n17 VP.n7 0.379447
R9971 VP.n356 VP.n355 0.379447
R9972 VP.n351 VP.n350 0.379447
R9973 VP.n346 VP.n345 0.379447
R9974 VP.n397 VP.n396 0.379447
R9975 VP.n392 VP.n391 0.379447
R9976 VP.n64 VP.n56 0.375125
R9977 VP.n85 VP.n49 0.375125
R9978 VP.n107 VP.n106 0.375125
R9979 VP.n126 VP.n122 0.375125
R9980 VP.n214 VP.n213 0.375125
R9981 VP.n291 VP.n229 0.375125
R9982 VP.n272 VP.n236 0.375125
R9983 VP.n249 VP.n246 0.375125
R9984 VP.n83 VP.n51 0.36275
R9985 VP.n100 VP.n45 0.36275
R9986 VP.n132 VP.n131 0.36275
R9987 VP.n297 VP.n296 0.36275
R9988 VP.n278 VP.n277 0.36275
R9989 VP.n254 VP.n244 0.36275
R9990 VP.n13 VP.n12 0.3605
R9991 VP.n19 VP.n18 0.3605
R9992 VP.n196 VP.n195 0.3605
R9993 VP.n189 VP.n28 0.3605
R9994 VP.n187 VP.n30 0.3605
R9995 VP.n177 VP.n33 0.3605
R9996 VP.n175 VP.n35 0.3605
R9997 VP.n170 VP.n38 0.3605
R9998 VP.n157 VP.n142 0.3605
R9999 VP.n152 VP.n145 0.3605
R10000 VP.n313 VP.n312 0.3605
R10001 VP.n319 VP.n318 0.3605
R10002 VP.n373 VP.n372 0.3605
R10003 VP.n366 VP.n328 0.3605
R10004 VP.n364 VP.n330 0.3605
R10005 VP.n354 VP.n333 0.3605
R10006 VP.n352 VP.n335 0.3605
R10007 VP.n347 VP.n338 0.3605
R10008 VP.n398 VP.n383 0.3605
R10009 VP.n393 VP.n386 0.3605
R10010 VP.n125 VP.n124 0.348488
R10011 VP.n248 VP.n247 0.348488
R10012 VP.n311 VP.n310 0.327481
R10013 VP.n11 VP.n10 0.327481
R10014 VP.n111 VP.n42 0.302474
R10015 VP.n93 VP.n48 0.302474
R10016 VP.n68 VP.n67 0.302474
R10017 VP.n269 VP.n268 0.302474
R10018 VP.n288 VP.n287 0.302474
R10019 VP.n218 VP.n206 0.302474
R10020 VP.n66 VP.n54 0.287375
R10021 VP.n92 VP.n91 0.287375
R10022 VP.n113 VP.n112 0.287375
R10023 VP.n220 VP.n219 0.287375
R10024 VP.n286 VP.n232 0.287375
R10025 VP.n267 VP.n239 0.287375
R10026 VP.n181 VP.n33 0.208099
R10027 VP.n358 VP.n333 0.208099
R10028 VP VP.n401 0.153263
R10029 VP.n377 VP.n376 0.147342
R10030 VP.n370 VP.n327 0.147342
R10031 VP.n367 VP.n329 0.147342
R10032 VP.n362 VP.n361 0.147342
R10033 VP.n315 VP.n314 0.147342
R10034 VP.n321 VP.n307 0.147342
R10035 VP.n134 VP.n133 0.147342
R10036 VP.n129 VP.n128 0.147342
R10037 VP.n101 VP.n46 0.147342
R10038 VP.n104 VP.n44 0.147342
R10039 VP.n111 VP.n110 0.147342
R10040 VP.n115 VP.n42 0.147342
R10041 VP.n80 VP.n79 0.147342
R10042 VP.n86 VP.n50 0.147342
R10043 VP.n89 VP.n48 0.147342
R10044 VP.n94 VP.n93 0.147342
R10045 VP.n61 VP.n60 0.147342
R10046 VP.n67 VP.n55 0.147342
R10047 VP.n69 VP.n68 0.147342
R10048 VP.n160 VP.n141 0.147342
R10049 VP.n155 VP.n154 0.147342
R10050 VP.n150 VP.n149 0.147342
R10051 VP.n178 VP.n34 0.147342
R10052 VP.n173 VP.n172 0.147342
R10053 VP.n168 VP.n167 0.147342
R10054 VP.n200 VP.n199 0.147342
R10055 VP.n193 VP.n27 0.147342
R10056 VP.n190 VP.n29 0.147342
R10057 VP.n185 VP.n184 0.147342
R10058 VP.n15 VP.n14 0.147342
R10059 VP.n21 VP.n7 0.147342
R10060 VP.n257 VP.n256 0.147342
R10061 VP.n252 VP.n251 0.147342
R10062 VP.n280 VP.n279 0.147342
R10063 VP.n275 VP.n274 0.147342
R10064 VP.n270 VP.n269 0.147342
R10065 VP.n268 VP.n240 0.147342
R10066 VP.n299 VP.n298 0.147342
R10067 VP.n294 VP.n293 0.147342
R10068 VP.n289 VP.n288 0.147342
R10069 VP.n287 VP.n233 0.147342
R10070 VP.n211 VP.n208 0.147342
R10071 VP.n218 VP.n217 0.147342
R10072 VP.n222 VP.n206 0.147342
R10073 VP.n355 VP.n334 0.147342
R10074 VP.n350 VP.n349 0.147342
R10075 VP.n345 VP.n344 0.147342
R10076 VP.n401 VP.n1 0.147342
R10077 VP.n396 VP.n395 0.147342
R10078 VP.n391 VP.n390 0.147342
R10079 VP.n375 VP.n374 0.142605
R10080 VP.n369 VP.n368 0.142605
R10081 VP.n363 VP.n331 0.142605
R10082 VP.n310 VP.n309 0.142605
R10083 VP.n317 VP.n316 0.142605
R10084 VP.n323 VP.n322 0.142605
R10085 VP.n156 VP.n143 0.142605
R10086 VP.n151 VP.n144 0.142605
R10087 VP.n180 VP.n179 0.142605
R10088 VP.n174 VP.n36 0.142605
R10089 VP.n169 VP.n37 0.142605
R10090 VP.n164 VP.n39 0.142605
R10091 VP.n198 VP.n197 0.142605
R10092 VP.n192 VP.n191 0.142605
R10093 VP.n186 VP.n31 0.142605
R10094 VP.n10 VP.n9 0.142605
R10095 VP.n17 VP.n16 0.142605
R10096 VP.n23 VP.n22 0.142605
R10097 VP.n357 VP.n356 0.142605
R10098 VP.n351 VP.n336 0.142605
R10099 VP.n346 VP.n337 0.142605
R10100 VP.n342 VP.n341 0.142605
R10101 VP.n397 VP.n384 0.142605
R10102 VP.n392 VP.n385 0.142605
R10103 VP.n59 VP.n56 0.14
R10104 VP.n65 VP.n64 0.14
R10105 VP.n66 VP.n65 0.14
R10106 VP.n70 VP.n54 0.14
R10107 VP.n71 VP.n70 0.14
R10108 VP.n78 VP.n77 0.14
R10109 VP.n78 VP.n51 0.14
R10110 VP.n84 VP.n83 0.14
R10111 VP.n85 VP.n84 0.14
R10112 VP.n90 VP.n49 0.14
R10113 VP.n91 VP.n90 0.14
R10114 VP.n92 VP.n47 0.14
R10115 VP.n96 VP.n47 0.14
R10116 VP.n99 VP.n98 0.14
R10117 VP.n100 VP.n99 0.14
R10118 VP.n105 VP.n45 0.14
R10119 VP.n106 VP.n105 0.14
R10120 VP.n107 VP.n43 0.14
R10121 VP.n112 VP.n43 0.14
R10122 VP.n114 VP.n113 0.14
R10123 VP.n114 VP.n40 0.14
R10124 VP.n137 VP.n41 0.14
R10125 VP.n132 VP.n41 0.14
R10126 VP.n131 VP.n130 0.14
R10127 VP.n130 VP.n122 0.14
R10128 VP.n13 VP.n8 0.14
R10129 VP.n18 VP.n8 0.14
R10130 VP.n20 VP.n19 0.14
R10131 VP.n20 VP.n5 0.14
R10132 VP.n201 VP.n6 0.14
R10133 VP.n196 VP.n6 0.14
R10134 VP.n195 VP.n194 0.14
R10135 VP.n194 VP.n28 0.14
R10136 VP.n189 VP.n188 0.14
R10137 VP.n188 VP.n187 0.14
R10138 VP.n183 VP.n30 0.14
R10139 VP.n183 VP.n182 0.14
R10140 VP.n177 VP.n176 0.14
R10141 VP.n176 VP.n175 0.14
R10142 VP.n171 VP.n35 0.14
R10143 VP.n171 VP.n170 0.14
R10144 VP.n166 VP.n38 0.14
R10145 VP.n166 VP.n165 0.14
R10146 VP.n159 VP.n158 0.14
R10147 VP.n158 VP.n157 0.14
R10148 VP.n153 VP.n142 0.14
R10149 VP.n153 VP.n152 0.14
R10150 VP.n148 VP.n145 0.14
R10151 VP.n213 VP.n212 0.14
R10152 VP.n214 VP.n207 0.14
R10153 VP.n219 VP.n207 0.14
R10154 VP.n221 VP.n220 0.14
R10155 VP.n221 VP.n204 0.14
R10156 VP.n302 VP.n205 0.14
R10157 VP.n297 VP.n205 0.14
R10158 VP.n296 VP.n295 0.14
R10159 VP.n295 VP.n229 0.14
R10160 VP.n291 VP.n290 0.14
R10161 VP.n290 VP.n232 0.14
R10162 VP.n286 VP.n285 0.14
R10163 VP.n285 VP.n284 0.14
R10164 VP.n282 VP.n234 0.14
R10165 VP.n278 VP.n234 0.14
R10166 VP.n277 VP.n276 0.14
R10167 VP.n276 VP.n236 0.14
R10168 VP.n272 VP.n271 0.14
R10169 VP.n271 VP.n239 0.14
R10170 VP.n267 VP.n266 0.14
R10171 VP.n266 VP.n265 0.14
R10172 VP.n259 VP.n258 0.14
R10173 VP.n258 VP.n244 0.14
R10174 VP.n254 VP.n253 0.14
R10175 VP.n253 VP.n246 0.14
R10176 VP.n313 VP.n308 0.14
R10177 VP.n318 VP.n308 0.14
R10178 VP.n320 VP.n319 0.14
R10179 VP.n320 VP.n305 0.14
R10180 VP.n378 VP.n306 0.14
R10181 VP.n373 VP.n306 0.14
R10182 VP.n372 VP.n371 0.14
R10183 VP.n371 VP.n328 0.14
R10184 VP.n366 VP.n365 0.14
R10185 VP.n365 VP.n364 0.14
R10186 VP.n360 VP.n330 0.14
R10187 VP.n360 VP.n359 0.14
R10188 VP.n354 VP.n353 0.14
R10189 VP.n353 VP.n352 0.14
R10190 VP.n348 VP.n335 0.14
R10191 VP.n348 VP.n347 0.14
R10192 VP.n343 VP.n338 0.14
R10193 VP.n343 VP.n2 0.14
R10194 VP.n400 VP.n399 0.14
R10195 VP.n399 VP.n398 0.14
R10196 VP.n394 VP.n383 0.14
R10197 VP.n394 VP.n393 0.14
R10198 VP.n389 VP.n386 0.14
R10199 VP.n117 VP.n116 0.118921
R10200 VP.n72 VP.n53 0.118921
R10201 VP.n264 VP.n242 0.118921
R10202 VP.n224 VP.n223 0.118921
R10203 VP.n136 VP.n135 0.116553
R10204 VP.n76 VP.n52 0.116553
R10205 VP.n260 VP.n243 0.116553
R10206 VP.n301 VP.n300 0.116553
R10207 VP.n123 VP.n121 0.114184
R10208 VP.n103 VP.n102 0.114184
R10209 VP.n82 VP.n81 0.114184
R10210 VP.n255 VP.n245 0.114184
R10211 VP.n237 VP.n235 0.114184
R10212 VP.n230 VP.n228 0.114184
R10213 VP.n127 VP.n124 0.0987895
R10214 VP.n109 VP.n108 0.0987895
R10215 VP.n88 VP.n87 0.0987895
R10216 VP.n63 VP.n62 0.0987895
R10217 VP.n250 VP.n247 0.0987895
R10218 VP.n273 VP.n238 0.0987895
R10219 VP.n292 VP.n231 0.0987895
R10220 VP.n216 VP.n215 0.0987895
R10221 VP.n110 VP.n109 0.0490526
R10222 VP.n89 VP.n88 0.0490526
R10223 VP.n62 VP.n55 0.0490526
R10224 VP.n270 VP.n238 0.0490526
R10225 VP.n289 VP.n231 0.0490526
R10226 VP.n217 VP.n216 0.0490526
R10227 VP.n129 VP.n123 0.0336579
R10228 VP.n104 VP.n103 0.0336579
R10229 VP.n81 VP.n50 0.0336579
R10230 VP.n60 VP.n57 0.0336579
R10231 VP.n252 VP.n245 0.0336579
R10232 VP.n275 VP.n237 0.0336579
R10233 VP.n294 VP.n230 0.0336579
R10234 VP.n211 VP.n210 0.0336579
R10235 VP.n135 VP.n134 0.0312895
R10236 VP.n97 VP.n46 0.0312895
R10237 VP.n79 VP.n52 0.0312895
R10238 VP.n257 VP.n243 0.0312895
R10239 VP.n281 VP.n280 0.0312895
R10240 VP.n300 VP.n299 0.0312895
R10241 VP.n116 VP.n115 0.0289211
R10242 VP.n95 VP.n94 0.0289211
R10243 VP.n69 VP.n53 0.0289211
R10244 VP.n242 VP.n240 0.0289211
R10245 VP.n283 VP.n233 0.0289211
R10246 VP.n223 VP.n222 0.0289211
R10247 VP.n376 VP.n375 0.00523684
R10248 VP.n370 VP.n369 0.00523684
R10249 VP.n331 VP.n329 0.00523684
R10250 VP.n361 VP.n332 0.00523684
R10251 VP.n316 VP.n315 0.00523684
R10252 VP.n322 VP.n321 0.00523684
R10253 VP.n143 VP.n141 0.00523684
R10254 VP.n154 VP.n144 0.00523684
R10255 VP.n149 VP.n146 0.00523684
R10256 VP.n36 VP.n34 0.00523684
R10257 VP.n172 VP.n37 0.00523684
R10258 VP.n167 VP.n39 0.00523684
R10259 VP.n199 VP.n198 0.00523684
R10260 VP.n193 VP.n192 0.00523684
R10261 VP.n31 VP.n29 0.00523684
R10262 VP.n184 VP.n32 0.00523684
R10263 VP.n16 VP.n15 0.00523684
R10264 VP.n22 VP.n21 0.00523684
R10265 VP.n336 VP.n334 0.00523684
R10266 VP.n349 VP.n337 0.00523684
R10267 VP.n344 VP.n342 0.00523684
R10268 VP.n384 VP.n1 0.00523684
R10269 VP.n395 VP.n385 0.00523684
R10270 VP.n390 VP.n387 0.00523684
R10271 a_n13990_n6451.n138 a_n13990_n6451.n137 8.18538
R10272 a_n13990_n6451.n62 a_n13990_n6451.n60 7.22198
R10273 a_n13990_n6451.n153 a_n13990_n6451.n152 7.22198
R10274 a_n13990_n6451.n47 a_n13990_n6451.t81 6.77653
R10275 a_n13990_n6451.n27 a_n13990_n6451.t56 6.77653
R10276 a_n13990_n6451.n82 a_n13990_n6451.t122 6.7761
R10277 a_n13990_n6451.n39 a_n13990_n6451.t134 6.7761
R10278 a_n13990_n6451.n25 a_n13990_n6451.t10 6.86989
R10279 a_n13990_n6451.n9 a_n13990_n6451.t116 6.77231
R10280 a_n13990_n6451.n19 a_n13990_n6451.t72 6.77231
R10281 a_n13990_n6451.n133 a_n13990_n6451.t36 6.53862
R10282 a_n13990_n6451.n145 a_n13990_n6451.n138 5.95467
R10283 a_n13990_n6451.n103 a_n13990_n6451.n101 5.89898
R10284 a_n13990_n6451.n117 a_n13990_n6451.t27 5.66511
R10285 a_n13990_n6451.n110 a_n13990_n6451.t50 5.66511
R10286 a_n13990_n6451.n118 a_n13990_n6451.t15 5.66379
R10287 a_n13990_n6451.n111 a_n13990_n6451.t1 5.66379
R10288 a_n13990_n6451.n110 a_n13990_n6451.n109 5.65285
R10289 a_n13990_n6451.n97 a_n13990_n6451.t5 5.61877
R10290 a_n13990_n6451.n98 a_n13990_n6451.t51 5.61877
R10291 a_n13990_n6451.n94 a_n13990_n6451.t8 5.61877
R10292 a_n13990_n6451.n79 a_n13990_n6451.t107 5.50607
R10293 a_n13990_n6451.n28 a_n13990_n6451.t85 5.50607
R10294 a_n13990_n6451.n51 a_n13990_n6451.t95 5.50607
R10295 a_n13990_n6451.n48 a_n13990_n6451.t130 5.50607
R10296 a_n13990_n6451.n80 a_n13990_n6451.t135 5.50475
R10297 a_n13990_n6451.n76 a_n13990_n6451.t89 5.50475
R10298 a_n13990_n6451.n75 a_n13990_n6451.t62 5.50475
R10299 a_n13990_n6451.n50 a_n13990_n6451.t58 5.50475
R10300 a_n13990_n6451.n54 a_n13990_n6451.t74 5.50475
R10301 a_n13990_n6451.n55 a_n13990_n6451.t77 5.50475
R10302 a_n13990_n6451.n49 a_n13990_n6451.t113 5.50475
R10303 a_n13990_n6451.t140 a_n13990_n6451.n157 5.50475
R10304 a_n13990_n6451.n136 a_n13990_n6451.t31 5.28484
R10305 a_n13990_n6451.n22 a_n13990_n6451.n123 5.29079
R10306 a_n13990_n6451.n120 a_n13990_n6451.n119 4.88835
R10307 a_n13990_n6451.n87 a_n13990_n6451.n86 4.88517
R10308 a_n13990_n6451.n124 a_n13990_n6451.n21 4.02009
R10309 a_n13990_n6451.t41 a_n13990_n6451.n20 5.28011
R10310 a_n13990_n6451.t46 a_n13990_n6451.n22 5.28011
R10311 a_n13990_n6451.n0 a_n13990_n6451.n72 4.0312
R10312 a_n13990_n6451.t93 a_n13990_n6451.n1 5.5012
R10313 a_n13990_n6451.t97 a_n13990_n6451.n2 5.5012
R10314 a_n13990_n6451.n71 a_n13990_n6451.n3 4.0312
R10315 a_n13990_n6451.t104 a_n13990_n6451.n4 5.5012
R10316 a_n13990_n6451.t114 a_n13990_n6451.n5 5.5012
R10317 a_n13990_n6451.n70 a_n13990_n6451.n6 4.0312
R10318 a_n13990_n6451.t55 a_n13990_n6451.n7 5.5012
R10319 a_n13990_n6451.t70 a_n13990_n6451.n8 5.5012
R10320 a_n13990_n6451.n68 a_n13990_n6451.n9 4.0312
R10321 a_n13990_n6451.n10 a_n13990_n6451.n143 4.0312
R10322 a_n13990_n6451.t60 a_n13990_n6451.n11 5.5012
R10323 a_n13990_n6451.t120 a_n13990_n6451.n12 5.5012
R10324 a_n13990_n6451.n142 a_n13990_n6451.n13 4.0312
R10325 a_n13990_n6451.t102 a_n13990_n6451.n14 5.5012
R10326 a_n13990_n6451.t76 a_n13990_n6451.n15 5.5012
R10327 a_n13990_n6451.n141 a_n13990_n6451.n16 4.0312
R10328 a_n13990_n6451.t67 a_n13990_n6451.n17 5.5012
R10329 a_n13990_n6451.t101 a_n13990_n6451.n18 5.5012
R10330 a_n13990_n6451.n139 a_n13990_n6451.n19 4.0312
R10331 a_n13990_n6451.n23 a_n13990_n6451.n96 4.40099
R10332 a_n13990_n6451.n24 a_n13990_n6451.n95 4.40099
R10333 a_n13990_n6451.n93 a_n13990_n6451.n25 4.40099
R10334 a_n13990_n6451.n116 a_n13990_n6451.n115 4.40379
R10335 a_n13990_n6451.n114 a_n13990_n6451.n113 4.40379
R10336 a_n13990_n6451.n102 a_n13990_n6451.t18 4.40142
R10337 a_n13990_n6451.n88 a_n13990_n6451.t11 4.40142
R10338 a_n13990_n6451.n61 a_n13990_n6451.t110 4.24002
R10339 a_n13990_n6451.n41 a_n13990_n6451.t82 4.24002
R10340 a_n13990_n6451.n151 a_n13990_n6451.t98 4.24002
R10341 a_n13990_n6451.n33 a_n13990_n6451.t103 4.24002
R10342 a_n13990_n6451.n129 a_n13990_n6451.t44 4.22616
R10343 a_n13990_n6451.n82 a_n13990_n6451.n81 4.03475
R10344 a_n13990_n6451.n78 a_n13990_n6451.n77 4.03475
R10345 a_n13990_n6451.n30 a_n13990_n6451.n29 4.03475
R10346 a_n13990_n6451.n27 a_n13990_n6451.n26 4.03475
R10347 a_n13990_n6451.n39 a_n13990_n6451.n38 4.03475
R10348 a_n13990_n6451.n53 a_n13990_n6451.n52 4.03475
R10349 a_n13990_n6451.n57 a_n13990_n6451.n56 4.03475
R10350 a_n13990_n6451.n47 a_n13990_n6451.n46 4.03475
R10351 a_n13990_n6451.n135 a_n13990_n6451.n134 4.02484
R10352 a_n13990_n6451.n133 a_n13990_n6451.n132 4.02484
R10353 a_n13990_n6451.n129 a_n13990_n6451.t38 4.02247
R10354 a_n13990_n6451.n131 a_n13990_n6451.n130 3.96014
R10355 a_n13990_n6451.n122 a_n13990_n6451.n85 3.94195
R10356 a_n13990_n6451.n102 a_n13990_n6451.t20 3.84721
R10357 a_n13990_n6451.n88 a_n13990_n6451.t4 3.84721
R10358 a_n13990_n6451.n116 a_n13990_n6451.n114 3.81703
R10359 a_n13990_n6451.n135 a_n13990_n6451.n133 3.80578
R10360 a_n13990_n6451.n61 a_n13990_n6451.t109 3.68818
R10361 a_n13990_n6451.n41 a_n13990_n6451.t80 3.68818
R10362 a_n13990_n6451.n151 a_n13990_n6451.t99 3.68818
R10363 a_n13990_n6451.n33 a_n13990_n6451.t105 3.68818
R10364 a_n13990_n6451.n67 a_n13990_n6451.n66 3.23904
R10365 a_n13990_n6451.n150 a_n13990_n6451.n146 3.23904
R10366 a_n13990_n6451.n108 a_n13990_n6451.n107 3.23004
R10367 a_n13990_n6451.n106 a_n13990_n6451.n105 3.14142
R10368 a_n13990_n6451.n91 a_n13990_n6451.n90 3.14142
R10369 a_n13990_n6451.n128 a_n13990_n6451.n126 2.96616
R10370 a_n13990_n6451.n65 a_n13990_n6451.n64 2.77002
R10371 a_n13990_n6451.n44 a_n13990_n6451.n43 2.77002
R10372 a_n13990_n6451.n149 a_n13990_n6451.n148 2.77002
R10373 a_n13990_n6451.n36 a_n13990_n6451.n35 2.77002
R10374 a_n13990_n6451.n128 a_n13990_n6451.n127 2.76247
R10375 a_n13990_n6451.n45 a_n13990_n6451.n41 2.73714
R10376 a_n13990_n6451.n37 a_n13990_n6451.n33 2.73714
R10377 a_n13990_n6451.n130 a_n13990_n6451.n128 2.71914
R10378 a_n13990_n6451.n92 a_n13990_n6451.n88 2.71914
R10379 a_n13990_n6451.n122 a_n13990_n6451.n121 2.64424
R10380 a_n13990_n6451.n55 a_n13990_n6451.n54 2.60203
R10381 a_n13990_n6451.n76 a_n13990_n6451.n75 2.60203
R10382 a_n13990_n6451.n106 a_n13990_n6451.n104 2.58721
R10383 a_n13990_n6451.n91 a_n13990_n6451.n89 2.58721
R10384 a_n13990_n6451.n111 a_n13990_n6451.n110 2.55136
R10385 a_n13990_n6451.n118 a_n13990_n6451.n117 2.55136
R10386 a_n13990_n6451.n157 a_n13990_n6451.n28 2.52471
R10387 a_n13990_n6451.n49 a_n13990_n6451.n48 2.52436
R10388 a_n13990_n6451.n51 a_n13990_n6451.n50 2.52436
R10389 a_n13990_n6451.n80 a_n13990_n6451.n79 2.52436
R10390 a_n13990_n6451.n100 a_n13990_n6451.n99 2.2807
R10391 a_n13990_n6451.n108 a_n13990_n6451.n87 2.2807
R10392 a_n13990_n6451.n65 a_n13990_n6451.n63 2.21818
R10393 a_n13990_n6451.n44 a_n13990_n6451.n42 2.21818
R10394 a_n13990_n6451.n149 a_n13990_n6451.n147 2.21818
R10395 a_n13990_n6451.n36 a_n13990_n6451.n34 2.21818
R10396 a_n13990_n6451.n59 a_n13990_n6451.n58 2.13841
R10397 a_n13990_n6451.n67 a_n13990_n6451.n40 2.13841
R10398 a_n13990_n6451.n60 a_n13990_n6451.n45 1.73904
R10399 a_n13990_n6451.n153 a_n13990_n6451.n37 1.73904
R10400 a_n13990_n6451.n137 a_n13990_n6451.n136 1.73609
R10401 a_n13990_n6451.n101 a_n13990_n6451.n92 1.73004
R10402 a_n13990_n6451.n140 a_n13990_n6451.n32 1.5005
R10403 a_n13990_n6451.n154 a_n13990_n6451.n153 1.5005
R10404 a_n13990_n6451.n69 a_n13990_n6451.n31 1.5005
R10405 a_n13990_n6451.n60 a_n13990_n6451.n59 1.5005
R10406 a_n13990_n6451.n101 a_n13990_n6451.n100 1.5005
R10407 a_n13990_n6451.n112 a_n13990_n6451.n85 1.5005
R10408 a_n13990_n6451.n121 a_n13990_n6451.n120 1.5005
R10409 a_n13990_n6451.n145 a_n13990_n6451.n144 1.5005
R10410 a_n13990_n6451.n74 a_n13990_n6451.n73 1.5005
R10411 a_n13990_n6451.n84 a_n13990_n6451.n83 1.5005
R10412 a_n13990_n6451.n156 a_n13990_n6451.n155 1.5005
R10413 a_n13990_n6451.n81 a_n13990_n6451.t66 1.4705
R10414 a_n13990_n6451.n81 a_n13990_n6451.t126 1.4705
R10415 a_n13990_n6451.n77 a_n13990_n6451.t115 1.4705
R10416 a_n13990_n6451.n77 a_n13990_n6451.t78 1.4705
R10417 a_n13990_n6451.n29 a_n13990_n6451.t71 1.4705
R10418 a_n13990_n6451.n29 a_n13990_n6451.t133 1.4705
R10419 a_n13990_n6451.n26 a_n13990_n6451.t108 1.4705
R10420 a_n13990_n6451.n26 a_n13990_n6451.t84 1.4705
R10421 a_n13990_n6451.n38 a_n13990_n6451.t65 1.4705
R10422 a_n13990_n6451.n38 a_n13990_n6451.t106 1.4705
R10423 a_n13990_n6451.n52 a_n13990_n6451.t137 1.4705
R10424 a_n13990_n6451.n52 a_n13990_n6451.t118 1.4705
R10425 a_n13990_n6451.n56 a_n13990_n6451.t119 1.4705
R10426 a_n13990_n6451.n56 a_n13990_n6451.t73 1.4705
R10427 a_n13990_n6451.n46 a_n13990_n6451.t75 1.4705
R10428 a_n13990_n6451.n46 a_n13990_n6451.t68 1.4705
R10429 a_n13990_n6451.n63 a_n13990_n6451.t139 1.4705
R10430 a_n13990_n6451.n63 a_n13990_n6451.t111 1.4705
R10431 a_n13990_n6451.n64 a_n13990_n6451.t141 1.4705
R10432 a_n13990_n6451.n64 a_n13990_n6451.t112 1.4705
R10433 a_n13990_n6451.n42 a_n13990_n6451.t86 1.4705
R10434 a_n13990_n6451.n42 a_n13990_n6451.t59 1.4705
R10435 a_n13990_n6451.n43 a_n13990_n6451.t88 1.4705
R10436 a_n13990_n6451.n43 a_n13990_n6451.t61 1.4705
R10437 a_n13990_n6451.n72 a_n13990_n6451.t129 1.4705
R10438 a_n13990_n6451.n72 a_n13990_n6451.t117 1.4705
R10439 a_n13990_n6451.n71 a_n13990_n6451.t69 1.4705
R10440 a_n13990_n6451.n71 a_n13990_n6451.t131 1.4705
R10441 a_n13990_n6451.n70 a_n13990_n6451.t91 1.4705
R10442 a_n13990_n6451.n70 a_n13990_n6451.t83 1.4705
R10443 a_n13990_n6451.n68 a_n13990_n6451.t90 1.4705
R10444 a_n13990_n6451.n68 a_n13990_n6451.t127 1.4705
R10445 a_n13990_n6451.n147 a_n13990_n6451.t96 1.4705
R10446 a_n13990_n6451.n147 a_n13990_n6451.t125 1.4705
R10447 a_n13990_n6451.n148 a_n13990_n6451.t94 1.4705
R10448 a_n13990_n6451.n148 a_n13990_n6451.t123 1.4705
R10449 a_n13990_n6451.n34 a_n13990_n6451.t124 1.4705
R10450 a_n13990_n6451.n34 a_n13990_n6451.t64 1.4705
R10451 a_n13990_n6451.n35 a_n13990_n6451.t121 1.4705
R10452 a_n13990_n6451.n35 a_n13990_n6451.t63 1.4705
R10453 a_n13990_n6451.n143 a_n13990_n6451.t79 1.4705
R10454 a_n13990_n6451.n143 a_n13990_n6451.t138 1.4705
R10455 a_n13990_n6451.n142 a_n13990_n6451.t132 1.4705
R10456 a_n13990_n6451.n142 a_n13990_n6451.t92 1.4705
R10457 a_n13990_n6451.n141 a_n13990_n6451.t87 1.4705
R10458 a_n13990_n6451.n141 a_n13990_n6451.t54 1.4705
R10459 a_n13990_n6451.n139 a_n13990_n6451.t128 1.4705
R10460 a_n13990_n6451.n139 a_n13990_n6451.t100 1.4705
R10461 a_n13990_n6451.n66 a_n13990_n6451.n65 1.46537
R10462 a_n13990_n6451.n62 a_n13990_n6451.n61 1.46537
R10463 a_n13990_n6451.n45 a_n13990_n6451.n44 1.46537
R10464 a_n13990_n6451.n150 a_n13990_n6451.n149 1.46537
R10465 a_n13990_n6451.n152 a_n13990_n6451.n151 1.46537
R10466 a_n13990_n6451.n37 a_n13990_n6451.n36 1.46537
R10467 a_n13990_n6451.n107 a_n13990_n6451.n106 1.46537
R10468 a_n13990_n6451.n103 a_n13990_n6451.n102 1.46537
R10469 a_n13990_n6451.n92 a_n13990_n6451.n91 1.46537
R10470 a_n13990_n6451.n130 a_n13990_n6451.n129 1.46537
R10471 a_n13990_n6451.n138 a_n13990_n6451.n32 1.37875
R10472 a_n13990_n6451.n57 a_n13990_n6451.n55 1.27228
R10473 a_n13990_n6451.n54 a_n13990_n6451.n53 1.27228
R10474 a_n13990_n6451.n66 a_n13990_n6451.n62 1.27228
R10475 a_n13990_n6451.n152 a_n13990_n6451.n150 1.27228
R10476 a_n13990_n6451.n75 a_n13990_n6451.n30 1.27228
R10477 a_n13990_n6451.n78 a_n13990_n6451.n76 1.27228
R10478 a_n13990_n6451.n48 a_n13990_n6451.n47 1.26756
R10479 a_n13990_n6451.n53 a_n13990_n6451.n51 1.26756
R10480 a_n13990_n6451.n28 a_n13990_n6451.n27 1.26756
R10481 a_n13990_n6451.n79 a_n13990_n6451.n78 1.26756
R10482 a_n13990_n6451.n125 a_n13990_n6451.n122 1.26344
R10483 a_n13990_n6451.n134 a_n13990_n6451.t32 1.2605
R10484 a_n13990_n6451.n134 a_n13990_n6451.t37 1.2605
R10485 a_n13990_n6451.n132 a_n13990_n6451.t40 1.2605
R10486 a_n13990_n6451.n132 a_n13990_n6451.t35 1.2605
R10487 a_n13990_n6451.n124 a_n13990_n6451.t42 1.2605
R10488 a_n13990_n6451.n124 a_n13990_n6451.t48 1.2605
R10489 a_n13990_n6451.n123 a_n13990_n6451.t47 1.2605
R10490 a_n13990_n6451.n123 a_n13990_n6451.t34 1.2605
R10491 a_n13990_n6451.n126 a_n13990_n6451.t45 1.2605
R10492 a_n13990_n6451.n126 a_n13990_n6451.t33 1.2605
R10493 a_n13990_n6451.n127 a_n13990_n6451.t39 1.2605
R10494 a_n13990_n6451.n127 a_n13990_n6451.t43 1.2605
R10495 a_n13990_n6451.n86 a_n13990_n6451.t26 1.2605
R10496 a_n13990_n6451.n86 a_n13990_n6451.t6 1.2605
R10497 a_n13990_n6451.n96 a_n13990_n6451.t7 1.2605
R10498 a_n13990_n6451.n96 a_n13990_n6451.t28 1.2605
R10499 a_n13990_n6451.n95 a_n13990_n6451.t30 1.2605
R10500 a_n13990_n6451.n95 a_n13990_n6451.t21 1.2605
R10501 a_n13990_n6451.n93 a_n13990_n6451.t25 1.2605
R10502 a_n13990_n6451.n93 a_n13990_n6451.t22 1.2605
R10503 a_n13990_n6451.n119 a_n13990_n6451.t23 1.2605
R10504 a_n13990_n6451.n119 a_n13990_n6451.t16 1.2605
R10505 a_n13990_n6451.n115 a_n13990_n6451.t14 1.2605
R10506 a_n13990_n6451.n115 a_n13990_n6451.t0 1.2605
R10507 a_n13990_n6451.n113 a_n13990_n6451.t19 1.2605
R10508 a_n13990_n6451.n113 a_n13990_n6451.t2 1.2605
R10509 a_n13990_n6451.n109 a_n13990_n6451.t29 1.2605
R10510 a_n13990_n6451.n109 a_n13990_n6451.t52 1.2605
R10511 a_n13990_n6451.n104 a_n13990_n6451.t13 1.2605
R10512 a_n13990_n6451.n104 a_n13990_n6451.t9 1.2605
R10513 a_n13990_n6451.n105 a_n13990_n6451.t53 1.2605
R10514 a_n13990_n6451.n105 a_n13990_n6451.t3 1.2605
R10515 a_n13990_n6451.n89 a_n13990_n6451.t24 1.2605
R10516 a_n13990_n6451.n89 a_n13990_n6451.t49 1.2605
R10517 a_n13990_n6451.n90 a_n13990_n6451.t17 1.2605
R10518 a_n13990_n6451.n90 a_n13990_n6451.t12 1.2605
R10519 a_n13990_n6451.n107 a_n13990_n6451.n103 1.25428
R10520 a_n13990_n6451.n136 a_n13990_n6451.n135 1.25428
R10521 a_n13990_n6451.n117 a_n13990_n6451.n116 1.24956
R10522 a_n13990_n6451.n98 a_n13990_n6451.n23 1.25162
R10523 a_n13990_n6451.n58 a_n13990_n6451.n49 0.796291
R10524 a_n13990_n6451.n50 a_n13990_n6451.n40 0.796291
R10525 a_n13990_n6451.n83 a_n13990_n6451.n80 0.796291
R10526 a_n13990_n6451.n157 a_n13990_n6451.n156 0.795934
R10527 a_n13990_n6451.n59 a_n13990_n6451.n31 0.780703
R10528 a_n13990_n6451.n154 a_n13990_n6451.n32 0.780703
R10529 a_n13990_n6451.n74 a_n13990_n6451.n67 0.780703
R10530 a_n13990_n6451.n146 a_n13990_n6451.n145 0.780703
R10531 a_n13990_n6451.n112 a_n13990_n6451.n111 0.769291
R10532 a_n13990_n6451.n120 a_n13990_n6451.n118 0.769291
R10533 a_n13990_n6451.n99 a_n13990_n6451.n94 0.767125
R10534 a_n13990_n6451.n97 a_n13990_n6451.n87 0.767125
R10535 a_n13990_n6451.n137 a_n13990_n6451.n131 0.639318
R10536 a_n13990_n6451.n155 a_n13990_n6451.n154 0.638405
R10537 a_n13990_n6451.n100 a_n13990_n6451.n85 0.638405
R10538 a_n13990_n6451.n121 a_n13990_n6451.n108 0.638405
R10539 a_n13990_n6451.n146 a_n13990_n6451.n84 0.638405
R10540 a_n13990_n6451.n155 a_n13990_n6451.n31 0.628372
R10541 a_n13990_n6451.n84 a_n13990_n6451.n74 0.628372
R10542 a_n13990_n6451.n131 a_n13990_n6451.n125 0.585196
R10543 a_n13990_n6451.n114 a_n13990_n6451.n112 0.485484
R10544 a_n13990_n6451.n58 a_n13990_n6451.n57 0.476484
R10545 a_n13990_n6451.n40 a_n13990_n6451.n39 0.476484
R10546 a_n13990_n6451.n156 a_n13990_n6451.n30 0.476484
R10547 a_n13990_n6451.n83 a_n13990_n6451.n82 0.476484
R10548 a_n13990_n6451.n99 a_n13990_n6451.n24 0.484998
R10549 a_n13990_n6451.n6 a_n13990_n6451.n69 0.478684
R10550 a_n13990_n6451.n73 a_n13990_n6451.n0 0.478684
R10551 a_n13990_n6451.n16 a_n13990_n6451.n140 0.478684
R10552 a_n13990_n6451.n144 a_n13990_n6451.n10 0.478684
R10553 a_n13990_n6451.n8 a_n13990_n6451.n9 1.27228
R10554 a_n13990_n6451.n7 a_n13990_n6451.n8 2.51878
R10555 a_n13990_n6451.n69 a_n13990_n6451.n7 0.794091
R10556 a_n13990_n6451.n5 a_n13990_n6451.n6 1.27228
R10557 a_n13990_n6451.n4 a_n13990_n6451.n5 2.60203
R10558 a_n13990_n6451.n3 a_n13990_n6451.n4 1.27228
R10559 a_n13990_n6451.n2 a_n13990_n6451.n3 1.27228
R10560 a_n13990_n6451.n1 a_n13990_n6451.n2 2.51878
R10561 a_n13990_n6451.n73 a_n13990_n6451.n1 0.794091
R10562 a_n13990_n6451.t57 a_n13990_n6451.n0 6.77266
R10563 a_n13990_n6451.n18 a_n13990_n6451.n19 1.27228
R10564 a_n13990_n6451.n17 a_n13990_n6451.n18 2.51878
R10565 a_n13990_n6451.n140 a_n13990_n6451.n17 0.794091
R10566 a_n13990_n6451.n15 a_n13990_n6451.n16 1.27228
R10567 a_n13990_n6451.n14 a_n13990_n6451.n15 2.60203
R10568 a_n13990_n6451.n13 a_n13990_n6451.n14 1.27228
R10569 a_n13990_n6451.n12 a_n13990_n6451.n13 1.27228
R10570 a_n13990_n6451.n11 a_n13990_n6451.n12 2.51878
R10571 a_n13990_n6451.n144 a_n13990_n6451.n11 0.794091
R10572 a_n13990_n6451.t136 a_n13990_n6451.n10 6.77266
R10573 a_n13990_n6451.n21 a_n13990_n6451.n22 3.15817
R10574 a_n13990_n6451.n20 a_n13990_n6451.n21 1.27188
R10575 a_n13990_n6451.n125 a_n13990_n6451.n20 1.73829
R10576 a_n13990_n6451.n94 a_n13990_n6451.n25 3.17898
R10577 a_n13990_n6451.n98 a_n13990_n6451.n24 3.19023
R10578 a_n13990_n6451.n97 a_n13990_n6451.n23 3.17898
R10579 VN.n0 VN.t28 8.10567
R10580 VN.n754 VN.t45 8.10567
R10581 VN.n36 VN.t12 8.10567
R10582 VN.n30 VN.t6 8.10567
R10583 VN.n49 VN.t62 8.10567
R10584 VN.n55 VN.t1 8.10567
R10585 VN.n786 VN.t67 8.10567
R10586 VN.n779 VN.t4 8.10567
R10587 VN.n835 VN.t58 8.10567
R10588 VN.n841 VN.t81 8.10567
R10589 VN.n190 VN.t21 8.10567
R10590 VN.n349 VN.t14 8.10567
R10591 VN.n343 VN.t38 8.10567
R10592 VN.n338 VN.t85 8.10567
R10593 VN.n333 VN.t2 8.10567
R10594 VN.n316 VN.t54 8.10567
R10595 VN.n305 VN.t31 8.10567
R10596 VN.n296 VN.t11 8.10567
R10597 VN.n287 VN.t72 8.10567
R10598 VN.n172 VN.t66 8.10567
R10599 VN.n267 VN.t75 8.10567
R10600 VN.n180 VN.t29 8.10567
R10601 VN.n184 VN.t34 8.10567
R10602 VN.n330 VN.t18 8.10567
R10603 VN.n323 VN.t80 8.10567
R10604 VN.n156 VN.t19 8.10567
R10605 VN.n246 VN.t69 8.10567
R10606 VN.n239 VN.t42 8.10567
R10607 VN.n188 VN.t51 8.10567
R10608 VN.n194 VN.t78 8.10567
R10609 VN.n212 VN.t70 8.10567
R10610 VN.n202 VN.t60 8.10567
R10611 VN.n100 VN.t20 8.10567
R10612 VN.n404 VN.t13 8.10567
R10613 VN.n398 VN.t37 8.10567
R10614 VN.n393 VN.t83 8.10567
R10615 VN.n389 VN.t0 8.10567
R10616 VN.n381 VN.t52 8.10567
R10617 VN.n144 VN.t30 8.10567
R10618 VN.n451 VN.t7 8.10567
R10619 VN.n457 VN.t71 8.10567
R10620 VN.n133 VN.t63 8.10567
R10621 VN.n126 VN.t73 8.10567
R10622 VN.n121 VN.t27 8.10567
R10623 VN.n478 VN.t33 8.10567
R10624 VN.n387 VN.t48 8.10567
R10625 VN.n386 VN.t17 8.10567
R10626 VN.n436 VN.t43 8.10567
R10627 VN.n114 VN.t82 8.10567
R10628 VN.n107 VN.t46 8.10567
R10629 VN.n65 VN.t84 8.10567
R10630 VN.n72 VN.t77 8.10567
R10631 VN.n74 VN.t68 8.10567
R10632 VN.n78 VN.t59 8.10567
R10633 VN.n532 VN.t44 8.10567
R10634 VN.n606 VN.t9 8.10567
R10635 VN.n600 VN.t5 8.10567
R10636 VN.n595 VN.t61 8.10567
R10637 VN.n590 VN.t87 8.10567
R10638 VN.n650 VN.t26 8.10567
R10639 VN.n660 VN.t55 8.10567
R10640 VN.n669 VN.t15 8.10567
R10641 VN.n678 VN.t40 8.10567
R10642 VN.n566 VN.t65 8.10567
R10643 VN.n559 VN.t3 8.10567
R10644 VN.n554 VN.t57 8.10567
R10645 VN.n549 VN.t79 8.10567
R10646 VN.n586 VN.t24 8.10567
R10647 VN.n585 VN.t53 8.10567
R10648 VN.n646 VN.t50 8.10567
R10649 VN.n546 VN.t86 8.10567
R10650 VN.n539 VN.t25 8.10567
R10651 VN.n489 VN.t39 8.10567
R10652 VN.n521 VN.t47 8.10567
R10653 VN.n512 VN.t22 8.10567
R10654 VN.n503 VN.t74 8.10567
R10655 VN.n743 VN.t49 8.10567
R10656 VN.n727 VN.t23 8.10567
R10657 VN.n730 VN.t76 8.10567
R10658 VN.n19 VN.t8 8.10567
R10659 VN.n12 VN.t36 8.10567
R10660 VN.n7 VN.t35 8.10567
R10661 VN.n768 VN.t64 8.10567
R10662 VN.n761 VN.t10 8.10567
R10663 VN.n719 VN.t32 8.10567
R10664 VN.n798 VN.t56 8.10567
R10665 VN.n793 VN.t16 8.10567
R10666 VN.n819 VN.t41 8.10567
R10667 VN.n846 VN.n845 7.83574
R10668 VN.n204 VN.n201 4.65575
R10669 VN.n505 VN.n502 4.65575
R10670 VN.n350 VN.n345 4.64641
R10671 VN.n607 VN.n604 4.64641
R10672 VN.n351 VN.n350 4.64
R10673 VN.n79 VN.n77 4.64
R10674 VN.n406 VN.n405 4.64
R10675 VN.n80 VN.n79 4.64
R10676 VN.n407 VN.n406 4.64
R10677 VN.n610 VN.n604 4.64
R10678 VN.n733 VN.n732 4.64
R10679 VN.n38 VN.n37 4.64
R10680 VN.n732 VN.n731 4.64
R10681 VN.n39 VN.n38 4.64
R10682 VN.n426 VN.n387 4.54125
R10683 VN.n115 VN.n114 4.54125
R10684 VN.n20 VN.n19 4.54125
R10685 VN.n769 VN.n768 4.54125
R10686 VN.n331 VN.n330 4.53893
R10687 VN.n247 VN.n246 4.53893
R10688 VN.n636 VN.n586 4.53893
R10689 VN.n547 VN.n546 4.53893
R10690 VN.n377 VN.n376 4.51011
R10691 VN.n284 VN.n170 4.51011
R10692 VN.n250 VN.n248 4.51011
R10693 VN.n634 VN.n589 4.51011
R10694 VN.n681 VN.n680 4.51011
R10695 VN.n711 VN.n710 4.51011
R10696 VN.n317 VN.n150 4.50691
R10697 VN.n283 VN.n282 4.50691
R10698 VN.n233 VN.n232 4.50691
R10699 VN.n649 VN.n580 4.50691
R10700 VN.n683 VN.n682 4.50691
R10701 VN.n533 VN.n483 4.50691
R10702 VN.n245 VN.n185 4.5005
R10703 VN.n244 VN.n243 4.5005
R10704 VN.n242 VN.n186 4.5005
R10705 VN.n241 VN.n240 4.5005
R10706 VN.n238 VN.n187 4.5005
R10707 VN.n237 VN.n236 4.5005
R10708 VN.n329 VN.n153 4.5005
R10709 VN.n328 VN.n327 4.5005
R10710 VN.n326 VN.n154 4.5005
R10711 VN.n325 VN.n324 4.5005
R10712 VN.n322 VN.n155 4.5005
R10713 VN.n321 VN.n320 4.5005
R10714 VN.n251 VN.n250 4.5005
R10715 VN.n253 VN.n252 4.5005
R10716 VN.n182 VN.n181 4.5005
R10717 VN.n260 VN.n259 4.5005
R10718 VN.n262 VN.n261 4.5005
R10719 VN.n178 VN.n177 4.5005
R10720 VN.n270 VN.n269 4.5005
R10721 VN.n271 VN.n176 4.5005
R10722 VN.n273 VN.n272 4.5005
R10723 VN.n174 VN.n173 4.5005
R10724 VN.n280 VN.n279 4.5005
R10725 VN.n282 VN.n281 4.5005
R10726 VN.n170 VN.n169 4.5005
R10727 VN.n289 VN.n288 4.5005
R10728 VN.n291 VN.n290 4.5005
R10729 VN.n166 VN.n165 4.5005
R10730 VN.n298 VN.n297 4.5005
R10731 VN.n300 VN.n299 4.5005
R10732 VN.n162 VN.n161 4.5005
R10733 VN.n308 VN.n307 4.5005
R10734 VN.n309 VN.n160 4.5005
R10735 VN.n311 VN.n310 4.5005
R10736 VN.n158 VN.n157 4.5005
R10737 VN.n318 VN.n317 4.5005
R10738 VN.n376 VN.n375 4.5005
R10739 VN.n374 VN.n373 4.5005
R10740 VN.n334 VN.n332 4.5005
R10741 VN.n368 VN.n367 4.5005
R10742 VN.n366 VN.n365 4.5005
R10743 VN.n339 VN.n337 4.5005
R10744 VN.n360 VN.n359 4.5005
R10745 VN.n358 VN.n357 4.5005
R10746 VN.n344 VN.n342 4.5005
R10747 VN.n348 VN.n346 4.5005
R10748 VN.n352 VN.n351 4.5005
R10749 VN.n204 VN.n203 4.5005
R10750 VN.n206 VN.n205 4.5005
R10751 VN.n198 VN.n197 4.5005
R10752 VN.n214 VN.n213 4.5005
R10753 VN.n216 VN.n215 4.5005
R10754 VN.n218 VN.n193 4.5005
R10755 VN.n224 VN.n223 4.5005
R10756 VN.n225 VN.n192 4.5005
R10757 VN.n227 VN.n226 4.5005
R10758 VN.n229 VN.n189 4.5005
R10759 VN.n234 VN.n233 4.5005
R10760 VN.n200 VN.n199 4.5005
R10761 VN.n208 VN.n207 4.5005
R10762 VN.n211 VN.n210 4.5005
R10763 VN.n209 VN.n196 4.5005
R10764 VN.n217 VN.n195 4.5005
R10765 VN.n220 VN.n219 4.5005
R10766 VN.n222 VN.n221 4.5005
R10767 VN.n228 VN.n191 4.5005
R10768 VN.n231 VN.n230 4.5005
R10769 VN.n249 VN.n183 4.5005
R10770 VN.n255 VN.n254 4.5005
R10771 VN.n257 VN.n256 4.5005
R10772 VN.n258 VN.n179 4.5005
R10773 VN.n264 VN.n263 4.5005
R10774 VN.n266 VN.n265 4.5005
R10775 VN.n268 VN.n175 4.5005
R10776 VN.n275 VN.n274 4.5005
R10777 VN.n277 VN.n276 4.5005
R10778 VN.n278 VN.n171 4.5005
R10779 VN.n286 VN.n285 4.5005
R10780 VN.n168 VN.n167 4.5005
R10781 VN.n293 VN.n292 4.5005
R10782 VN.n295 VN.n294 4.5005
R10783 VN.n164 VN.n163 4.5005
R10784 VN.n302 VN.n301 4.5005
R10785 VN.n304 VN.n303 4.5005
R10786 VN.n306 VN.n159 4.5005
R10787 VN.n313 VN.n312 4.5005
R10788 VN.n315 VN.n314 4.5005
R10789 VN.n152 VN.n151 4.5005
R10790 VN.n372 VN.n371 4.5005
R10791 VN.n370 VN.n369 4.5005
R10792 VN.n336 VN.n335 4.5005
R10793 VN.n364 VN.n363 4.5005
R10794 VN.n362 VN.n361 4.5005
R10795 VN.n341 VN.n340 4.5005
R10796 VN.n356 VN.n355 4.5005
R10797 VN.n354 VN.n353 4.5005
R10798 VN.n347 VN.n345 4.5005
R10799 VN.n113 VN.n62 4.5005
R10800 VN.n112 VN.n111 4.5005
R10801 VN.n110 VN.n63 4.5005
R10802 VN.n109 VN.n108 4.5005
R10803 VN.n106 VN.n64 4.5005
R10804 VN.n105 VN.n104 4.5005
R10805 VN.n428 VN.n427 4.5005
R10806 VN.n429 VN.n385 4.5005
R10807 VN.n431 VN.n430 4.5005
R10808 VN.n432 VN.n384 4.5005
R10809 VN.n434 VN.n433 4.5005
R10810 VN.n435 VN.n383 4.5005
R10811 VN.n461 VN.n460 4.5005
R10812 VN.n134 VN.n131 4.5005
R10813 VN.n465 VN.n130 4.5005
R10814 VN.n466 VN.n129 4.5005
R10815 VN.n467 VN.n128 4.5005
R10816 VN.n470 VN.n125 4.5005
R10817 VN.n471 VN.n124 4.5005
R10818 VN.n472 VN.n123 4.5005
R10819 VN.n122 VN.n119 4.5005
R10820 VN.n476 VN.n118 4.5005
R10821 VN.n477 VN.n117 4.5005
R10822 VN.n479 VN.n116 4.5005
R10823 VN.n439 VN.n438 4.5005
R10824 VN.n382 VN.n149 4.5005
R10825 VN.n443 VN.n148 4.5005
R10826 VN.n444 VN.n147 4.5005
R10827 VN.n445 VN.n146 4.5005
R10828 VN.n145 VN.n142 4.5005
R10829 VN.n449 VN.n141 4.5005
R10830 VN.n450 VN.n140 4.5005
R10831 VN.n452 VN.n139 4.5005
R10832 VN.n138 VN.n136 4.5005
R10833 VN.n456 VN.n135 4.5005
R10834 VN.n459 VN.n458 4.5005
R10835 VN.n405 VN.n403 4.5005
R10836 VN.n409 VN.n402 4.5005
R10837 VN.n410 VN.n401 4.5005
R10838 VN.n411 VN.n400 4.5005
R10839 VN.n414 VN.n397 4.5005
R10840 VN.n415 VN.n396 4.5005
R10841 VN.n416 VN.n395 4.5005
R10842 VN.n419 VN.n392 4.5005
R10843 VN.n420 VN.n391 4.5005
R10844 VN.n421 VN.n388 4.5005
R10845 VN.n425 VN.n424 4.5005
R10846 VN.n102 VN.n101 4.5005
R10847 VN.n99 VN.n66 4.5005
R10848 VN.n93 VN.n67 4.5005
R10849 VN.n95 VN.n94 4.5005
R10850 VN.n92 VN.n69 4.5005
R10851 VN.n91 VN.n90 4.5005
R10852 VN.n71 VN.n70 4.5005
R10853 VN.n86 VN.n85 4.5005
R10854 VN.n84 VN.n83 4.5005
R10855 VN.n82 VN.n75 4.5005
R10856 VN.n77 VN.n76 4.5005
R10857 VN.n80 VN.n76 4.5005
R10858 VN.n82 VN.n81 4.5005
R10859 VN.n83 VN.n73 4.5005
R10860 VN.n87 VN.n86 4.5005
R10861 VN.n88 VN.n71 4.5005
R10862 VN.n90 VN.n89 4.5005
R10863 VN.n69 VN.n68 4.5005
R10864 VN.n96 VN.n95 4.5005
R10865 VN.n97 VN.n67 4.5005
R10866 VN.n99 VN.n98 4.5005
R10867 VN.n101 VN.n60 4.5005
R10868 VN.n480 VN.n479 4.5005
R10869 VN.n477 VN.n61 4.5005
R10870 VN.n476 VN.n475 4.5005
R10871 VN.n474 VN.n119 4.5005
R10872 VN.n473 VN.n472 4.5005
R10873 VN.n471 VN.n120 4.5005
R10874 VN.n470 VN.n469 4.5005
R10875 VN.n468 VN.n467 4.5005
R10876 VN.n466 VN.n127 4.5005
R10877 VN.n465 VN.n464 4.5005
R10878 VN.n463 VN.n131 4.5005
R10879 VN.n462 VN.n461 4.5005
R10880 VN.n458 VN.n132 4.5005
R10881 VN.n456 VN.n455 4.5005
R10882 VN.n454 VN.n136 4.5005
R10883 VN.n453 VN.n452 4.5005
R10884 VN.n450 VN.n137 4.5005
R10885 VN.n449 VN.n448 4.5005
R10886 VN.n447 VN.n142 4.5005
R10887 VN.n446 VN.n445 4.5005
R10888 VN.n444 VN.n143 4.5005
R10889 VN.n443 VN.n442 4.5005
R10890 VN.n441 VN.n149 4.5005
R10891 VN.n440 VN.n439 4.5005
R10892 VN.n424 VN.n423 4.5005
R10893 VN.n422 VN.n421 4.5005
R10894 VN.n420 VN.n390 4.5005
R10895 VN.n419 VN.n418 4.5005
R10896 VN.n417 VN.n416 4.5005
R10897 VN.n415 VN.n394 4.5005
R10898 VN.n414 VN.n413 4.5005
R10899 VN.n412 VN.n411 4.5005
R10900 VN.n410 VN.n399 4.5005
R10901 VN.n409 VN.n408 4.5005
R10902 VN.n407 VN.n403 4.5005
R10903 VN.n545 VN.n486 4.5005
R10904 VN.n544 VN.n543 4.5005
R10905 VN.n542 VN.n487 4.5005
R10906 VN.n541 VN.n540 4.5005
R10907 VN.n538 VN.n488 4.5005
R10908 VN.n537 VN.n536 4.5005
R10909 VN.n638 VN.n637 4.5005
R10910 VN.n639 VN.n584 4.5005
R10911 VN.n641 VN.n640 4.5005
R10912 VN.n642 VN.n583 4.5005
R10913 VN.n644 VN.n643 4.5005
R10914 VN.n645 VN.n582 4.5005
R10915 VN.n710 VN.n709 4.5005
R10916 VN.n708 VN.n707 4.5005
R10917 VN.n550 VN.n548 4.5005
R10918 VN.n702 VN.n701 4.5005
R10919 VN.n700 VN.n699 4.5005
R10920 VN.n555 VN.n553 4.5005
R10921 VN.n694 VN.n693 4.5005
R10922 VN.n692 VN.n691 4.5005
R10923 VN.n560 VN.n558 4.5005
R10924 VN.n564 VN.n562 4.5005
R10925 VN.n686 VN.n685 4.5005
R10926 VN.n684 VN.n683 4.5005
R10927 VN.n680 VN.n565 4.5005
R10928 VN.n677 VN.n676 4.5005
R10929 VN.n675 VN.n674 4.5005
R10930 VN.n570 VN.n569 4.5005
R10931 VN.n668 VN.n667 4.5005
R10932 VN.n666 VN.n665 4.5005
R10933 VN.n575 VN.n574 4.5005
R10934 VN.n659 VN.n658 4.5005
R10935 VN.n657 VN.n656 4.5005
R10936 VN.n655 VN.n578 4.5005
R10937 VN.n581 VN.n579 4.5005
R10938 VN.n649 VN.n648 4.5005
R10939 VN.n635 VN.n634 4.5005
R10940 VN.n592 VN.n587 4.5005
R10941 VN.n629 VN.n628 4.5005
R10942 VN.n627 VN.n626 4.5005
R10943 VN.n597 VN.n594 4.5005
R10944 VN.n621 VN.n620 4.5005
R10945 VN.n619 VN.n618 4.5005
R10946 VN.n602 VN.n599 4.5005
R10947 VN.n613 VN.n612 4.5005
R10948 VN.n611 VN.n603 4.5005
R10949 VN.n610 VN.n609 4.5005
R10950 VN.n505 VN.n504 4.5005
R10951 VN.n507 VN.n506 4.5005
R10952 VN.n499 VN.n498 4.5005
R10953 VN.n514 VN.n513 4.5005
R10954 VN.n516 VN.n515 4.5005
R10955 VN.n495 VN.n494 4.5005
R10956 VN.n524 VN.n523 4.5005
R10957 VN.n525 VN.n493 4.5005
R10958 VN.n527 VN.n526 4.5005
R10959 VN.n491 VN.n490 4.5005
R10960 VN.n534 VN.n533 4.5005
R10961 VN.n501 VN.n500 4.5005
R10962 VN.n509 VN.n508 4.5005
R10963 VN.n511 VN.n510 4.5005
R10964 VN.n497 VN.n496 4.5005
R10965 VN.n518 VN.n517 4.5005
R10966 VN.n520 VN.n519 4.5005
R10967 VN.n522 VN.n492 4.5005
R10968 VN.n529 VN.n528 4.5005
R10969 VN.n531 VN.n530 4.5005
R10970 VN.n485 VN.n484 4.5005
R10971 VN.n706 VN.n705 4.5005
R10972 VN.n704 VN.n703 4.5005
R10973 VN.n552 VN.n551 4.5005
R10974 VN.n698 VN.n697 4.5005
R10975 VN.n696 VN.n695 4.5005
R10976 VN.n557 VN.n556 4.5005
R10977 VN.n690 VN.n689 4.5005
R10978 VN.n688 VN.n687 4.5005
R10979 VN.n563 VN.n561 4.5005
R10980 VN.n679 VN.n567 4.5005
R10981 VN.n571 VN.n568 4.5005
R10982 VN.n673 VN.n672 4.5005
R10983 VN.n671 VN.n670 4.5005
R10984 VN.n573 VN.n572 4.5005
R10985 VN.n664 VN.n663 4.5005
R10986 VN.n662 VN.n661 4.5005
R10987 VN.n577 VN.n576 4.5005
R10988 VN.n654 VN.n653 4.5005
R10989 VN.n652 VN.n651 4.5005
R10990 VN.n633 VN.n632 4.5005
R10991 VN.n631 VN.n630 4.5005
R10992 VN.n593 VN.n591 4.5005
R10993 VN.n625 VN.n624 4.5005
R10994 VN.n623 VN.n622 4.5005
R10995 VN.n598 VN.n596 4.5005
R10996 VN.n617 VN.n616 4.5005
R10997 VN.n615 VN.n614 4.5005
R10998 VN.n605 VN.n601 4.5005
R10999 VN.n608 VN.n607 4.5005
R11000 VN.n843 VN.n842 4.5005
R11001 VN.n840 VN.n715 4.5005
R11002 VN.n773 VN.n771 4.5005
R11003 VN.n836 VN.n774 4.5005
R11004 VN.n834 VN.n775 4.5005
R11005 VN.n833 VN.n776 4.5005
R11006 VN.n780 VN.n777 4.5005
R11007 VN.n829 VN.n781 4.5005
R11008 VN.n828 VN.n782 4.5005
R11009 VN.n827 VN.n783 4.5005
R11010 VN.n787 VN.n784 4.5005
R11011 VN.n823 VN.n822 4.5005
R11012 VN.n57 VN.n56 4.5005
R11013 VN.n54 VN.n3 4.5005
R11014 VN.n24 VN.n22 4.5005
R11015 VN.n50 VN.n25 4.5005
R11016 VN.n48 VN.n26 4.5005
R11017 VN.n47 VN.n27 4.5005
R11018 VN.n31 VN.n28 4.5005
R11019 VN.n43 VN.n32 4.5005
R11020 VN.n42 VN.n33 4.5005
R11021 VN.n41 VN.n34 4.5005
R11022 VN.n37 VN.n35 4.5005
R11023 VN.n733 VN.n729 4.5005
R11024 VN.n735 VN.n734 4.5005
R11025 VN.n736 VN.n726 4.5005
R11026 VN.n740 VN.n739 4.5005
R11027 VN.n741 VN.n725 4.5005
R11028 VN.n744 VN.n742 4.5005
R11029 VN.n723 VN.n722 4.5005
R11030 VN.n750 VN.n749 4.5005
R11031 VN.n751 VN.n721 4.5005
R11032 VN.n753 VN.n752 4.5005
R11033 VN.n755 VN.n714 4.5005
R11034 VN.n767 VN.n716 4.5005
R11035 VN.n766 VN.n765 4.5005
R11036 VN.n764 VN.n717 4.5005
R11037 VN.n763 VN.n762 4.5005
R11038 VN.n760 VN.n718 4.5005
R11039 VN.n759 VN.n758 4.5005
R11040 VN.n18 VN.n4 4.5005
R11041 VN.n17 VN.n16 4.5005
R11042 VN.n15 VN.n5 4.5005
R11043 VN.n14 VN.n13 4.5005
R11044 VN.n11 VN.n6 4.5005
R11045 VN.n10 VN.n9 4.5005
R11046 VN.n756 VN.n755 4.5005
R11047 VN.n753 VN.n720 4.5005
R11048 VN.n747 VN.n721 4.5005
R11049 VN.n749 VN.n748 4.5005
R11050 VN.n746 VN.n723 4.5005
R11051 VN.n745 VN.n744 4.5005
R11052 VN.n725 VN.n724 4.5005
R11053 VN.n739 VN.n738 4.5005
R11054 VN.n737 VN.n736 4.5005
R11055 VN.n735 VN.n728 4.5005
R11056 VN.n731 VN.n729 4.5005
R11057 VN.n824 VN.n823 4.5005
R11058 VN.n825 VN.n784 4.5005
R11059 VN.n827 VN.n826 4.5005
R11060 VN.n828 VN.n778 4.5005
R11061 VN.n830 VN.n829 4.5005
R11062 VN.n831 VN.n777 4.5005
R11063 VN.n833 VN.n832 4.5005
R11064 VN.n834 VN.n772 4.5005
R11065 VN.n837 VN.n836 4.5005
R11066 VN.n838 VN.n771 4.5005
R11067 VN.n840 VN.n839 4.5005
R11068 VN.n842 VN.n770 4.5005
R11069 VN.n39 VN.n35 4.5005
R11070 VN.n41 VN.n40 4.5005
R11071 VN.n42 VN.n29 4.5005
R11072 VN.n44 VN.n43 4.5005
R11073 VN.n45 VN.n28 4.5005
R11074 VN.n47 VN.n46 4.5005
R11075 VN.n48 VN.n23 4.5005
R11076 VN.n51 VN.n50 4.5005
R11077 VN.n52 VN.n22 4.5005
R11078 VN.n54 VN.n53 4.5005
R11079 VN.n56 VN.n21 4.5005
R11080 VN.n849 VN.n1 4.5005
R11081 VN.n804 VN.n803 4.5005
R11082 VN.n806 VN.n802 4.5005
R11083 VN.n807 VN.n801 4.5005
R11084 VN.n808 VN.n800 4.5005
R11085 VN.n811 VN.n797 4.5005
R11086 VN.n812 VN.n796 4.5005
R11087 VN.n813 VN.n795 4.5005
R11088 VN.n794 VN.n791 4.5005
R11089 VN.n817 VN.n790 4.5005
R11090 VN.n818 VN.n789 4.5005
R11091 VN.n820 VN.n785 4.5005
R11092 VN.n821 VN.n820 4.5005
R11093 VN.n818 VN.n788 4.5005
R11094 VN.n817 VN.n816 4.5005
R11095 VN.n815 VN.n791 4.5005
R11096 VN.n814 VN.n813 4.5005
R11097 VN.n812 VN.n792 4.5005
R11098 VN.n811 VN.n810 4.5005
R11099 VN.n809 VN.n808 4.5005
R11100 VN.n807 VN.n799 4.5005
R11101 VN.n806 VN.n805 4.5005
R11102 VN.n804 VN.n2 4.5005
R11103 VN.n849 VN.n848 4.5005
R11104 VN.n281 VN.n169 3.0245
R11105 VN.n460 VN.n459 3.0245
R11106 VN.n462 VN.n132 3.0245
R11107 VN.n684 VN.n565 3.0245
R11108 VN.n822 VN.n821 3.0245
R11109 VN.n824 VN.n785 3.0245
R11110 VN.n284 VN.n283 2.96825
R11111 VN.n682 VN.n681 2.96825
R11112 VN.n201 VN.n199 2.41967
R11113 VN.n502 VN.n500 2.41967
R11114 VN.n437 VN.n436 2.22849
R11115 VN.n103 VN.n65 2.22849
R11116 VN.n8 VN.n7 2.22849
R11117 VN.n757 VN.n719 2.22849
R11118 VN.n319 VN.n156 2.22782
R11119 VN.n235 VN.n188 2.22782
R11120 VN.n647 VN.n646 2.22782
R11121 VN.n535 VN.n489 2.22782
R11122 VN.n481 VN.n480 2.102
R11123 VN.n423 VN.n380 2.102
R11124 VN.n844 VN.n843 2.102
R11125 VN.n847 VN.n57 2.102
R11126 VN.n482 VN.n59 2.07182
R11127 VN.n379 VN.n378 2.07182
R11128 VN.n248 VN.n59 2.06825
R11129 VN.n378 VN.n377 2.06825
R11130 VN.n712 VN.n711 2.06825
R11131 VN.n589 VN.n588 2.06825
R11132 VN.n713 VN.n712 1.5005
R11133 VN.n482 VN.n481 1.5005
R11134 VN.n588 VN.n58 1.5005
R11135 VN.n380 VN.n379 1.5005
R11136 VN.n847 VN.n846 1.5005
R11137 VN.n845 VN.n844 1.5005
R11138 VN.n713 VN.n482 1.47516
R11139 VN.n379 VN.n58 1.47516
R11140 VN.n481 VN.n60 0.83975
R11141 VN.n440 VN.n380 0.83975
R11142 VN.n844 VN.n714 0.83975
R11143 VN.n848 VN.n847 0.83975
R11144 VN.n232 VN.n59 0.81725
R11145 VN.n378 VN.n150 0.81725
R11146 VN.n712 VN.n483 0.81725
R11147 VN.n588 VN.n580 0.81725
R11148 VN.n103 VN.n102 0.75626
R11149 VN.n438 VN.n437 0.75626
R11150 VN.n757 VN.n756 0.75626
R11151 VN.n8 VN.n1 0.75626
R11152 VN.n235 VN.n234 0.756242
R11153 VN.n319 VN.n318 0.756242
R11154 VN.n535 VN.n534 0.756242
R11155 VN.n648 VN.n647 0.756242
R11156 VN.n251 VN.n247 0.698
R11157 VN.n375 VN.n331 0.698
R11158 VN.n116 VN.n115 0.698
R11159 VN.n426 VN.n425 0.698
R11160 VN.n709 VN.n547 0.698
R11161 VN.n636 VN.n635 0.698
R11162 VN.n770 VN.n769 0.698
R11163 VN.n21 VN.n20 0.698
R11164 VN.n845 VN.n713 0.571818
R11165 VN.n846 VN.n58 0.571818
R11166 VN.n215 VN.n193 0.375125
R11167 VN.n270 VN.n177 0.375125
R11168 VN.n299 VN.n161 0.375125
R11169 VN.n359 VN.n337 0.375125
R11170 VN.n91 VN.n70 0.375125
R11171 VN.n125 VN.n124 0.375125
R11172 VN.n145 VN.n141 0.375125
R11173 VN.n397 VN.n396 0.375125
R11174 VN.n89 VN.n88 0.375125
R11175 VN.n469 VN.n120 0.375125
R11176 VN.n448 VN.n447 0.375125
R11177 VN.n413 VN.n394 0.375125
R11178 VN.n515 VN.n494 0.375125
R11179 VN.n693 VN.n553 0.375125
R11180 VN.n666 VN.n574 0.375125
R11181 VN.n620 VN.n619 0.375125
R11182 VN.n742 VN.n741 0.375125
R11183 VN.n780 VN.n776 0.375125
R11184 VN.n810 VN.n792 0.375125
R11185 VN.n31 VN.n27 0.375125
R11186 VN.n745 VN.n724 0.375125
R11187 VN.n832 VN.n831 0.375125
R11188 VN.n797 VN.n796 0.375125
R11189 VN.n46 VN.n45 0.375125
R11190 VN.n205 VN.n197 0.36275
R11191 VN.n260 VN.n181 0.36275
R11192 VN.n290 VN.n165 0.36275
R11193 VN.n367 VN.n332 0.36275
R11194 VN.n84 VN.n75 0.36275
R11195 VN.n122 VN.n118 0.36275
R11196 VN.n139 VN.n138 0.36275
R11197 VN.n392 VN.n391 0.36275
R11198 VN.n81 VN.n73 0.36275
R11199 VN.n475 VN.n474 0.36275
R11200 VN.n454 VN.n453 0.36275
R11201 VN.n418 VN.n390 0.36275
R11202 VN.n506 VN.n498 0.36275
R11203 VN.n701 VN.n548 0.36275
R11204 VN.n675 VN.n569 0.36275
R11205 VN.n628 VN.n627 0.36275
R11206 VN.n734 VN.n726 0.36275
R11207 VN.n774 VN.n773 0.36275
R11208 VN.n816 VN.n815 0.36275
R11209 VN.n25 VN.n24 0.36275
R11210 VN.n737 VN.n728 0.36275
R11211 VN.n838 VN.n837 0.36275
R11212 VN.n794 VN.n790 0.36275
R11213 VN.n52 VN.n51 0.36275
R11214 VN.n236 VN.n187 0.3605
R11215 VN.n243 VN.n242 0.3605
R11216 VN.n320 VN.n155 0.3605
R11217 VN.n327 VN.n326 0.3605
R11218 VN.n208 VN.n199 0.3605
R11219 VN.n209 VN.n195 0.3605
R11220 VN.n221 VN.n191 0.3605
R11221 VN.n256 VN.n255 0.3605
R11222 VN.n265 VN.n264 0.3605
R11223 VN.n276 VN.n275 0.3605
R11224 VN.n293 VN.n167 0.3605
R11225 VN.n302 VN.n163 0.3605
R11226 VN.n313 VN.n159 0.3605
R11227 VN.n371 VN.n370 0.3605
R11228 VN.n363 VN.n362 0.3605
R11229 VN.n355 VN.n354 0.3605
R11230 VN.n104 VN.n64 0.3605
R11231 VN.n111 VN.n110 0.3605
R11232 VN.n433 VN.n383 0.3605
R11233 VN.n431 VN.n385 0.3605
R11234 VN.n536 VN.n488 0.3605
R11235 VN.n543 VN.n542 0.3605
R11236 VN.n643 VN.n582 0.3605
R11237 VN.n641 VN.n584 0.3605
R11238 VN.n509 VN.n500 0.3605
R11239 VN.n518 VN.n496 0.3605
R11240 VN.n529 VN.n492 0.3605
R11241 VN.n705 VN.n704 0.3605
R11242 VN.n697 VN.n696 0.3605
R11243 VN.n689 VN.n688 0.3605
R11244 VN.n672 VN.n571 0.3605
R11245 VN.n663 VN.n572 0.3605
R11246 VN.n653 VN.n576 0.3605
R11247 VN.n631 VN.n591 0.3605
R11248 VN.n623 VN.n596 0.3605
R11249 VN.n615 VN.n601 0.3605
R11250 VN.n758 VN.n718 0.3605
R11251 VN.n765 VN.n764 0.3605
R11252 VN.n9 VN.n6 0.3605
R11253 VN.n16 VN.n15 0.3605
R11254 VN.n226 VN.n225 0.287375
R11255 VN.n272 VN.n173 0.287375
R11256 VN.n310 VN.n309 0.287375
R11257 VN.n348 VN.n342 0.287375
R11258 VN.n94 VN.n93 0.287375
R11259 VN.n130 VN.n129 0.287375
R11260 VN.n148 VN.n147 0.287375
R11261 VN.n402 VN.n401 0.287375
R11262 VN.n97 VN.n96 0.287375
R11263 VN.n464 VN.n127 0.287375
R11264 VN.n442 VN.n143 0.287375
R11265 VN.n408 VN.n399 0.287375
R11266 VN.n526 VN.n525 0.287375
R11267 VN.n564 VN.n558 0.287375
R11268 VN.n657 VN.n578 0.287375
R11269 VN.n612 VN.n611 0.287375
R11270 VN.n751 VN.n750 0.287375
R11271 VN.n783 VN.n782 0.287375
R11272 VN.n805 VN.n799 0.287375
R11273 VN.n34 VN.n33 0.287375
R11274 VN.n748 VN.n747 0.287375
R11275 VN.n826 VN.n778 0.287375
R11276 VN.n802 VN.n801 0.287375
R11277 VN.n40 VN.n29 0.287375
R11278 VN.n236 VN.n235 0.208888
R11279 VN.n320 VN.n319 0.208888
R11280 VN.n536 VN.n535 0.208888
R11281 VN.n647 VN.n582 0.208888
R11282 VN.n104 VN.n103 0.20887
R11283 VN.n437 VN.n383 0.20887
R11284 VN.n758 VN.n757 0.20887
R11285 VN.n9 VN.n8 0.20887
R11286 VN.n205 VN.n204 0.14
R11287 VN.n214 VN.n197 0.14
R11288 VN.n215 VN.n214 0.14
R11289 VN.n224 VN.n193 0.14
R11290 VN.n225 VN.n224 0.14
R11291 VN.n226 VN.n189 0.14
R11292 VN.n234 VN.n189 0.14
R11293 VN.n241 VN.n187 0.14
R11294 VN.n242 VN.n241 0.14
R11295 VN.n243 VN.n185 0.14
R11296 VN.n247 VN.n185 0.14
R11297 VN.n252 VN.n251 0.14
R11298 VN.n252 VN.n181 0.14
R11299 VN.n261 VN.n260 0.14
R11300 VN.n261 VN.n177 0.14
R11301 VN.n271 VN.n270 0.14
R11302 VN.n272 VN.n271 0.14
R11303 VN.n280 VN.n173 0.14
R11304 VN.n281 VN.n280 0.14
R11305 VN.n289 VN.n169 0.14
R11306 VN.n290 VN.n289 0.14
R11307 VN.n298 VN.n165 0.14
R11308 VN.n299 VN.n298 0.14
R11309 VN.n308 VN.n161 0.14
R11310 VN.n309 VN.n308 0.14
R11311 VN.n310 VN.n157 0.14
R11312 VN.n318 VN.n157 0.14
R11313 VN.n325 VN.n155 0.14
R11314 VN.n326 VN.n325 0.14
R11315 VN.n327 VN.n153 0.14
R11316 VN.n331 VN.n153 0.14
R11317 VN.n375 VN.n374 0.14
R11318 VN.n374 VN.n332 0.14
R11319 VN.n367 VN.n366 0.14
R11320 VN.n366 VN.n337 0.14
R11321 VN.n359 VN.n358 0.14
R11322 VN.n358 VN.n342 0.14
R11323 VN.n351 VN.n348 0.14
R11324 VN.n210 VN.n208 0.14
R11325 VN.n210 VN.n209 0.14
R11326 VN.n220 VN.n195 0.14
R11327 VN.n221 VN.n220 0.14
R11328 VN.n231 VN.n191 0.14
R11329 VN.n232 VN.n231 0.14
R11330 VN.n248 VN.n183 0.14
R11331 VN.n255 VN.n183 0.14
R11332 VN.n256 VN.n179 0.14
R11333 VN.n264 VN.n179 0.14
R11334 VN.n265 VN.n175 0.14
R11335 VN.n275 VN.n175 0.14
R11336 VN.n276 VN.n171 0.14
R11337 VN.n283 VN.n171 0.14
R11338 VN.n285 VN.n284 0.14
R11339 VN.n285 VN.n167 0.14
R11340 VN.n294 VN.n293 0.14
R11341 VN.n294 VN.n163 0.14
R11342 VN.n303 VN.n302 0.14
R11343 VN.n303 VN.n159 0.14
R11344 VN.n314 VN.n313 0.14
R11345 VN.n314 VN.n150 0.14
R11346 VN.n377 VN.n151 0.14
R11347 VN.n371 VN.n151 0.14
R11348 VN.n370 VN.n335 0.14
R11349 VN.n363 VN.n335 0.14
R11350 VN.n362 VN.n340 0.14
R11351 VN.n355 VN.n340 0.14
R11352 VN.n354 VN.n345 0.14
R11353 VN.n77 VN.n75 0.14
R11354 VN.n85 VN.n84 0.14
R11355 VN.n85 VN.n70 0.14
R11356 VN.n92 VN.n91 0.14
R11357 VN.n94 VN.n92 0.14
R11358 VN.n93 VN.n66 0.14
R11359 VN.n102 VN.n66 0.14
R11360 VN.n109 VN.n64 0.14
R11361 VN.n110 VN.n109 0.14
R11362 VN.n111 VN.n62 0.14
R11363 VN.n115 VN.n62 0.14
R11364 VN.n117 VN.n116 0.14
R11365 VN.n118 VN.n117 0.14
R11366 VN.n123 VN.n122 0.14
R11367 VN.n124 VN.n123 0.14
R11368 VN.n128 VN.n125 0.14
R11369 VN.n129 VN.n128 0.14
R11370 VN.n134 VN.n130 0.14
R11371 VN.n460 VN.n134 0.14
R11372 VN.n459 VN.n135 0.14
R11373 VN.n138 VN.n135 0.14
R11374 VN.n140 VN.n139 0.14
R11375 VN.n141 VN.n140 0.14
R11376 VN.n146 VN.n145 0.14
R11377 VN.n147 VN.n146 0.14
R11378 VN.n382 VN.n148 0.14
R11379 VN.n438 VN.n382 0.14
R11380 VN.n433 VN.n432 0.14
R11381 VN.n432 VN.n431 0.14
R11382 VN.n427 VN.n385 0.14
R11383 VN.n427 VN.n426 0.14
R11384 VN.n425 VN.n388 0.14
R11385 VN.n391 VN.n388 0.14
R11386 VN.n395 VN.n392 0.14
R11387 VN.n396 VN.n395 0.14
R11388 VN.n400 VN.n397 0.14
R11389 VN.n401 VN.n400 0.14
R11390 VN.n405 VN.n402 0.14
R11391 VN.n81 VN.n80 0.14
R11392 VN.n87 VN.n73 0.14
R11393 VN.n88 VN.n87 0.14
R11394 VN.n89 VN.n68 0.14
R11395 VN.n96 VN.n68 0.14
R11396 VN.n98 VN.n97 0.14
R11397 VN.n98 VN.n60 0.14
R11398 VN.n480 VN.n61 0.14
R11399 VN.n475 VN.n61 0.14
R11400 VN.n474 VN.n473 0.14
R11401 VN.n473 VN.n120 0.14
R11402 VN.n469 VN.n468 0.14
R11403 VN.n468 VN.n127 0.14
R11404 VN.n464 VN.n463 0.14
R11405 VN.n463 VN.n462 0.14
R11406 VN.n455 VN.n132 0.14
R11407 VN.n455 VN.n454 0.14
R11408 VN.n453 VN.n137 0.14
R11409 VN.n448 VN.n137 0.14
R11410 VN.n447 VN.n446 0.14
R11411 VN.n446 VN.n143 0.14
R11412 VN.n442 VN.n441 0.14
R11413 VN.n441 VN.n440 0.14
R11414 VN.n423 VN.n422 0.14
R11415 VN.n422 VN.n390 0.14
R11416 VN.n418 VN.n417 0.14
R11417 VN.n417 VN.n394 0.14
R11418 VN.n413 VN.n412 0.14
R11419 VN.n412 VN.n399 0.14
R11420 VN.n408 VN.n407 0.14
R11421 VN.n506 VN.n505 0.14
R11422 VN.n514 VN.n498 0.14
R11423 VN.n515 VN.n514 0.14
R11424 VN.n524 VN.n494 0.14
R11425 VN.n525 VN.n524 0.14
R11426 VN.n526 VN.n490 0.14
R11427 VN.n534 VN.n490 0.14
R11428 VN.n541 VN.n488 0.14
R11429 VN.n542 VN.n541 0.14
R11430 VN.n543 VN.n486 0.14
R11431 VN.n547 VN.n486 0.14
R11432 VN.n709 VN.n708 0.14
R11433 VN.n708 VN.n548 0.14
R11434 VN.n701 VN.n700 0.14
R11435 VN.n700 VN.n553 0.14
R11436 VN.n693 VN.n692 0.14
R11437 VN.n692 VN.n558 0.14
R11438 VN.n685 VN.n564 0.14
R11439 VN.n685 VN.n684 0.14
R11440 VN.n676 VN.n565 0.14
R11441 VN.n676 VN.n675 0.14
R11442 VN.n667 VN.n569 0.14
R11443 VN.n667 VN.n666 0.14
R11444 VN.n658 VN.n574 0.14
R11445 VN.n658 VN.n657 0.14
R11446 VN.n581 VN.n578 0.14
R11447 VN.n648 VN.n581 0.14
R11448 VN.n643 VN.n642 0.14
R11449 VN.n642 VN.n641 0.14
R11450 VN.n637 VN.n584 0.14
R11451 VN.n637 VN.n636 0.14
R11452 VN.n635 VN.n587 0.14
R11453 VN.n628 VN.n587 0.14
R11454 VN.n627 VN.n594 0.14
R11455 VN.n620 VN.n594 0.14
R11456 VN.n619 VN.n599 0.14
R11457 VN.n612 VN.n599 0.14
R11458 VN.n611 VN.n610 0.14
R11459 VN.n510 VN.n509 0.14
R11460 VN.n510 VN.n496 0.14
R11461 VN.n519 VN.n518 0.14
R11462 VN.n519 VN.n492 0.14
R11463 VN.n530 VN.n529 0.14
R11464 VN.n530 VN.n483 0.14
R11465 VN.n711 VN.n484 0.14
R11466 VN.n705 VN.n484 0.14
R11467 VN.n704 VN.n551 0.14
R11468 VN.n697 VN.n551 0.14
R11469 VN.n696 VN.n556 0.14
R11470 VN.n689 VN.n556 0.14
R11471 VN.n688 VN.n561 0.14
R11472 VN.n682 VN.n561 0.14
R11473 VN.n681 VN.n567 0.14
R11474 VN.n571 VN.n567 0.14
R11475 VN.n672 VN.n671 0.14
R11476 VN.n671 VN.n572 0.14
R11477 VN.n663 VN.n662 0.14
R11478 VN.n662 VN.n576 0.14
R11479 VN.n653 VN.n652 0.14
R11480 VN.n652 VN.n580 0.14
R11481 VN.n632 VN.n589 0.14
R11482 VN.n632 VN.n631 0.14
R11483 VN.n624 VN.n591 0.14
R11484 VN.n624 VN.n623 0.14
R11485 VN.n616 VN.n596 0.14
R11486 VN.n616 VN.n615 0.14
R11487 VN.n607 VN.n601 0.14
R11488 VN.n734 VN.n733 0.14
R11489 VN.n740 VN.n726 0.14
R11490 VN.n741 VN.n740 0.14
R11491 VN.n742 VN.n722 0.14
R11492 VN.n750 VN.n722 0.14
R11493 VN.n752 VN.n751 0.14
R11494 VN.n752 VN.n714 0.14
R11495 VN.n843 VN.n715 0.14
R11496 VN.n773 VN.n715 0.14
R11497 VN.n775 VN.n774 0.14
R11498 VN.n776 VN.n775 0.14
R11499 VN.n781 VN.n780 0.14
R11500 VN.n782 VN.n781 0.14
R11501 VN.n787 VN.n783 0.14
R11502 VN.n822 VN.n787 0.14
R11503 VN.n821 VN.n788 0.14
R11504 VN.n816 VN.n788 0.14
R11505 VN.n815 VN.n814 0.14
R11506 VN.n814 VN.n792 0.14
R11507 VN.n810 VN.n809 0.14
R11508 VN.n809 VN.n799 0.14
R11509 VN.n805 VN.n2 0.14
R11510 VN.n848 VN.n2 0.14
R11511 VN.n57 VN.n3 0.14
R11512 VN.n24 VN.n3 0.14
R11513 VN.n26 VN.n25 0.14
R11514 VN.n27 VN.n26 0.14
R11515 VN.n32 VN.n31 0.14
R11516 VN.n33 VN.n32 0.14
R11517 VN.n37 VN.n34 0.14
R11518 VN.n731 VN.n728 0.14
R11519 VN.n738 VN.n737 0.14
R11520 VN.n738 VN.n724 0.14
R11521 VN.n746 VN.n745 0.14
R11522 VN.n748 VN.n746 0.14
R11523 VN.n747 VN.n720 0.14
R11524 VN.n756 VN.n720 0.14
R11525 VN.n763 VN.n718 0.14
R11526 VN.n764 VN.n763 0.14
R11527 VN.n765 VN.n716 0.14
R11528 VN.n769 VN.n716 0.14
R11529 VN.n839 VN.n770 0.14
R11530 VN.n839 VN.n838 0.14
R11531 VN.n837 VN.n772 0.14
R11532 VN.n832 VN.n772 0.14
R11533 VN.n831 VN.n830 0.14
R11534 VN.n830 VN.n778 0.14
R11535 VN.n826 VN.n825 0.14
R11536 VN.n825 VN.n824 0.14
R11537 VN.n789 VN.n785 0.14
R11538 VN.n790 VN.n789 0.14
R11539 VN.n795 VN.n794 0.14
R11540 VN.n796 VN.n795 0.14
R11541 VN.n800 VN.n797 0.14
R11542 VN.n801 VN.n800 0.14
R11543 VN.n803 VN.n802 0.14
R11544 VN.n803 VN.n1 0.14
R11545 VN.n14 VN.n6 0.14
R11546 VN.n15 VN.n14 0.14
R11547 VN.n16 VN.n4 0.14
R11548 VN.n20 VN.n4 0.14
R11549 VN.n53 VN.n21 0.14
R11550 VN.n53 VN.n52 0.14
R11551 VN.n51 VN.n23 0.14
R11552 VN.n46 VN.n23 0.14
R11553 VN.n45 VN.n44 0.14
R11554 VN.n44 VN.n29 0.14
R11555 VN.n40 VN.n39 0.14
R11556 VN.n435 VN.n434 0.109179
R11557 VN.n430 VN.n429 0.109179
R11558 VN.n106 VN.n105 0.109179
R11559 VN.n112 VN.n63 0.109179
R11560 VN.n11 VN.n10 0.109179
R11561 VN.n17 VN.n5 0.109179
R11562 VN.n760 VN.n759 0.109179
R11563 VN.n766 VN.n717 0.109179
R11564 VN.n47 VN.n28 0.107155
R11565 VN.n833 VN.n777 0.107155
R11566 VN.n415 VN.n414 0.107155
R11567 VN.n449 VN.n142 0.107155
R11568 VN.n471 VN.n470 0.107155
R11569 VN.n90 VN.n71 0.107155
R11570 VN.n744 VN.n725 0.107155
R11571 VN.n812 VN.n811 0.107155
R11572 VN.n50 VN.n22 0.103632
R11573 VN.n836 VN.n771 0.103632
R11574 VN.n420 VN.n419 0.103632
R11575 VN.n452 VN.n136 0.103632
R11576 VN.n476 VN.n119 0.103632
R11577 VN.n83 VN.n82 0.103632
R11578 VN.n736 VN.n735 0.103632
R11579 VN.n817 VN.n791 0.103632
R11580 VN.n322 VN.n321 0.102991
R11581 VN.n328 VN.n154 0.102991
R11582 VN.n238 VN.n237 0.102991
R11583 VN.n244 VN.n186 0.102991
R11584 VN.n645 VN.n644 0.102991
R11585 VN.n640 VN.n639 0.102991
R11586 VN.n538 VN.n537 0.102991
R11587 VN.n544 VN.n487 0.102991
R11588 VN.n369 VN.n334 0.0933826
R11589 VN.n292 VN.n291 0.0933826
R11590 VN.n257 VN.n182 0.0933826
R11591 VN.n207 VN.n206 0.0933826
R11592 VN.n629 VN.n593 0.0933826
R11593 VN.n674 VN.n673 0.0933826
R11594 VN.n703 VN.n550 0.0933826
R11595 VN.n508 VN.n507 0.0933826
R11596 VN.n361 VN.n339 0.092742
R11597 VN.n301 VN.n300 0.092742
R11598 VN.n266 VN.n178 0.092742
R11599 VN.n217 VN.n216 0.092742
R11600 VN.n621 VN.n598 0.092742
R11601 VN.n665 VN.n664 0.092742
R11602 VN.n695 VN.n555 0.092742
R11603 VN.n517 VN.n516 0.092742
R11604 VN.n42 VN.n41 0.0821726
R11605 VN.n828 VN.n827 0.0821726
R11606 VN.n346 VN.n344 0.0821726
R11607 VN.n311 VN.n160 0.0821726
R11608 VN.n273 VN.n174 0.0821726
R11609 VN.n227 VN.n192 0.0821726
R11610 VN.n410 VN.n409 0.0821726
R11611 VN.n444 VN.n443 0.0821726
R11612 VN.n466 VN.n465 0.0821726
R11613 VN.n95 VN.n67 0.0821726
R11614 VN.n613 VN.n603 0.0821726
R11615 VN.n656 VN.n655 0.0821726
R11616 VN.n562 VN.n560 0.0821726
R11617 VN.n527 VN.n493 0.0821726
R11618 VN.n749 VN.n721 0.0821726
R11619 VN.n807 VN.n806 0.0821726
R11620 VN.n434 VN.n384 0.0426132
R11621 VN.n429 VN.n428 0.0426132
R11622 VN.n108 VN.n106 0.0426132
R11623 VN.n113 VN.n112 0.0426132
R11624 VN.n13 VN.n11 0.0426132
R11625 VN.n18 VN.n17 0.0426132
R11626 VN.n762 VN.n760 0.0426132
R11627 VN.n767 VN.n766 0.0426132
R11628 VN.n436 VN.n435 0.0412547
R11629 VN.n430 VN.n386 0.0412547
R11630 VN.n105 VN.n65 0.0412547
R11631 VN.n107 VN.n63 0.0412547
R11632 VN.n10 VN.n7 0.0412547
R11633 VN.n12 VN.n5 0.0412547
R11634 VN.n759 VN.n719 0.0412547
R11635 VN.n761 VN.n717 0.0412547
R11636 VN.n54 VN.n22 0.0402153
R11637 VN.n48 VN.n47 0.0402153
R11638 VN.n43 VN.n42 0.0402153
R11639 VN.n41 VN.n35 0.0402153
R11640 VN.n840 VN.n771 0.0402153
R11641 VN.n834 VN.n833 0.0402153
R11642 VN.n829 VN.n828 0.0402153
R11643 VN.n827 VN.n784 0.0402153
R11644 VN.n324 VN.n322 0.0402153
R11645 VN.n329 VN.n328 0.0402153
R11646 VN.n240 VN.n238 0.0402153
R11647 VN.n245 VN.n244 0.0402153
R11648 VN.n421 VN.n420 0.0402153
R11649 VN.n416 VN.n415 0.0402153
R11650 VN.n411 VN.n410 0.0402153
R11651 VN.n409 VN.n403 0.0402153
R11652 VN.n456 VN.n136 0.0402153
R11653 VN.n450 VN.n449 0.0402153
R11654 VN.n445 VN.n444 0.0402153
R11655 VN.n443 VN.n149 0.0402153
R11656 VN.n477 VN.n476 0.0402153
R11657 VN.n472 VN.n471 0.0402153
R11658 VN.n467 VN.n466 0.0402153
R11659 VN.n465 VN.n131 0.0402153
R11660 VN.n82 VN.n76 0.0402153
R11661 VN.n86 VN.n71 0.0402153
R11662 VN.n95 VN.n69 0.0402153
R11663 VN.n99 VN.n67 0.0402153
R11664 VN.n644 VN.n583 0.0402153
R11665 VN.n639 VN.n638 0.0402153
R11666 VN.n540 VN.n538 0.0402153
R11667 VN.n545 VN.n544 0.0402153
R11668 VN.n735 VN.n729 0.0402153
R11669 VN.n739 VN.n725 0.0402153
R11670 VN.n749 VN.n723 0.0402153
R11671 VN.n753 VN.n721 0.0402153
R11672 VN.n818 VN.n817 0.0402153
R11673 VN.n813 VN.n812 0.0402153
R11674 VN.n808 VN.n807 0.0402153
R11675 VN.n806 VN.n804 0.0402153
R11676 VN.n321 VN.n156 0.0389342
R11677 VN.n323 VN.n154 0.0389342
R11678 VN.n237 VN.n188 0.0389342
R11679 VN.n239 VN.n186 0.0389342
R11680 VN.n646 VN.n645 0.0389342
R11681 VN.n640 VN.n585 0.0389342
R11682 VN.n537 VN.n489 0.0389342
R11683 VN.n539 VN.n487 0.0389342
R11684 VN.n353 VN.n352 0.0338096
R11685 VN.n312 VN.n158 0.0338096
R11686 VN.n279 VN.n277 0.0338096
R11687 VN.n229 VN.n228 0.0338096
R11688 VN.n609 VN.n605 0.0338096
R11689 VN.n654 VN.n579 0.0338096
R11690 VN.n687 VN.n686 0.0338096
R11691 VN.n528 VN.n491 0.0338096
R11692 VN.n38 VN.n36 0.0325285
R11693 VN.n823 VN.n786 0.0325285
R11694 VN.n350 VN.n349 0.0325285
R11695 VN.n317 VN.n316 0.0325285
R11696 VN.n282 VN.n172 0.0325285
R11697 VN.n233 VN.n190 0.0325285
R11698 VN.n406 VN.n404 0.0325285
R11699 VN.n439 VN.n381 0.0325285
R11700 VN.n461 VN.n133 0.0325285
R11701 VN.n101 VN.n100 0.0325285
R11702 VN.n606 VN.n604 0.0325285
R11703 VN.n650 VN.n649 0.0325285
R11704 VN.n683 VN.n566 0.0325285
R11705 VN.n533 VN.n532 0.0325285
R11706 VN.n755 VN.n754 0.0325285
R11707 VN.n849 VN.n0 0.0325285
R11708 VN.n56 VN.n55 0.0318879
R11709 VN.n842 VN.n841 0.0318879
R11710 VN.n424 VN.n389 0.0318879
R11711 VN.n458 VN.n457 0.0318879
R11712 VN.n479 VN.n478 0.0318879
R11713 VN.n79 VN.n78 0.0318879
R11714 VN.n732 VN.n730 0.0318879
R11715 VN.n820 VN.n819 0.0318879
R11716 VN.n50 VN.n49 0.0312473
R11717 VN.n836 VN.n835 0.0312473
R11718 VN.n419 VN.n393 0.0312473
R11719 VN.n452 VN.n451 0.0312473
R11720 VN.n121 VN.n119 0.0312473
R11721 VN.n83 VN.n74 0.0312473
R11722 VN.n736 VN.n727 0.0312473
R11723 VN.n793 VN.n791 0.0312473
R11724 VN.n376 VN.n152 0.0306068
R11725 VN.n373 VN.n372 0.0306068
R11726 VN.n286 VN.n170 0.0306068
R11727 VN.n288 VN.n168 0.0306068
R11728 VN.n250 VN.n249 0.0306068
R11729 VN.n254 VN.n253 0.0306068
R11730 VN.n203 VN.n200 0.0306068
R11731 VN.n634 VN.n633 0.0306068
R11732 VN.n630 VN.n592 0.0306068
R11733 VN.n680 VN.n679 0.0306068
R11734 VN.n677 VN.n568 0.0306068
R11735 VN.n710 VN.n485 0.0306068
R11736 VN.n707 VN.n706 0.0306068
R11737 VN.n504 VN.n501 0.0306068
R11738 VN.n368 VN.n336 0.0299662
R11739 VN.n365 VN.n364 0.0299662
R11740 VN.n295 VN.n166 0.0299662
R11741 VN.n297 VN.n164 0.0299662
R11742 VN.n259 VN.n258 0.0299662
R11743 VN.n263 VN.n262 0.0299662
R11744 VN.n211 VN.n198 0.0299662
R11745 VN.n213 VN.n196 0.0299662
R11746 VN.n626 VN.n625 0.0299662
R11747 VN.n622 VN.n597 0.0299662
R11748 VN.n670 VN.n570 0.0299662
R11749 VN.n668 VN.n573 0.0299662
R11750 VN.n702 VN.n552 0.0299662
R11751 VN.n699 VN.n698 0.0299662
R11752 VN.n511 VN.n499 0.0299662
R11753 VN.n513 VN.n497 0.0299662
R11754 VN.n30 VN.n28 0.0270836
R11755 VN.n779 VN.n777 0.0270836
R11756 VN.n414 VN.n398 0.0270836
R11757 VN.n144 VN.n142 0.0270836
R11758 VN.n470 VN.n126 0.0270836
R11759 VN.n90 VN.n72 0.0270836
R11760 VN.n744 VN.n743 0.0270836
R11761 VN.n811 VN.n798 0.0270836
R11762 VN.n360 VN.n341 0.0258025
R11763 VN.n357 VN.n356 0.0258025
R11764 VN.n304 VN.n162 0.0258025
R11765 VN.n307 VN.n306 0.0258025
R11766 VN.n269 VN.n268 0.0258025
R11767 VN.n274 VN.n176 0.0258025
R11768 VN.n219 VN.n218 0.0258025
R11769 VN.n223 VN.n222 0.0258025
R11770 VN.n618 VN.n617 0.0258025
R11771 VN.n614 VN.n602 0.0258025
R11772 VN.n661 VN.n575 0.0258025
R11773 VN.n659 VN.n577 0.0258025
R11774 VN.n694 VN.n557 0.0258025
R11775 VN.n691 VN.n690 0.0258025
R11776 VN.n520 VN.n495 0.0258025
R11777 VN.n523 VN.n522 0.0258025
R11778 VN.n202 VN.n201 0.0170406
R11779 VN.n503 VN.n502 0.0170406
R11780 VN.n361 VN.n360 0.0149128
R11781 VN.n356 VN.n344 0.0149128
R11782 VN.n301 VN.n162 0.0149128
R11783 VN.n306 VN.n160 0.0149128
R11784 VN.n269 VN.n266 0.0149128
R11785 VN.n274 VN.n273 0.0149128
R11786 VN.n218 VN.n217 0.0149128
R11787 VN.n222 VN.n192 0.0149128
R11788 VN.n618 VN.n598 0.0149128
R11789 VN.n614 VN.n613 0.0149128
R11790 VN.n664 VN.n575 0.0149128
R11791 VN.n656 VN.n577 0.0149128
R11792 VN.n695 VN.n694 0.0149128
R11793 VN.n690 VN.n560 0.0149128
R11794 VN.n517 VN.n495 0.0149128
R11795 VN.n522 VN.n493 0.0149128
R11796 VN.n43 VN.n30 0.0136317
R11797 VN.n829 VN.n779 0.0136317
R11798 VN.n357 VN.n343 0.0136317
R11799 VN.n307 VN.n305 0.0136317
R11800 VN.n267 VN.n176 0.0136317
R11801 VN.n223 VN.n194 0.0136317
R11802 VN.n411 VN.n398 0.0136317
R11803 VN.n445 VN.n144 0.0136317
R11804 VN.n467 VN.n126 0.0136317
R11805 VN.n72 VN.n69 0.0136317
R11806 VN.n602 VN.n600 0.0136317
R11807 VN.n660 VN.n659 0.0136317
R11808 VN.n691 VN.n559 0.0136317
R11809 VN.n523 VN.n521 0.0136317
R11810 VN.n743 VN.n723 0.0136317
R11811 VN.n808 VN.n798 0.0136317
R11812 VN.n369 VN.n368 0.0107491
R11813 VN.n364 VN.n339 0.0107491
R11814 VN.n292 VN.n166 0.0107491
R11815 VN.n300 VN.n164 0.0107491
R11816 VN.n259 VN.n257 0.0107491
R11817 VN.n263 VN.n178 0.0107491
R11818 VN.n207 VN.n198 0.0107491
R11819 VN.n216 VN.n196 0.0107491
R11820 VN.n626 VN.n593 0.0107491
R11821 VN.n622 VN.n621 0.0107491
R11822 VN.n673 VN.n570 0.0107491
R11823 VN.n665 VN.n573 0.0107491
R11824 VN.n703 VN.n702 0.0107491
R11825 VN.n698 VN.n555 0.0107491
R11826 VN.n508 VN.n499 0.0107491
R11827 VN.n516 VN.n497 0.0107491
R11828 VN.n372 VN.n334 0.0101085
R11829 VN.n291 VN.n168 0.0101085
R11830 VN.n254 VN.n182 0.0101085
R11831 VN.n206 VN.n200 0.0101085
R11832 VN.n630 VN.n629 0.0101085
R11833 VN.n674 VN.n568 0.0101085
R11834 VN.n706 VN.n550 0.0101085
R11835 VN.n507 VN.n501 0.0101085
R11836 VN.n49 VN.n48 0.00946797
R11837 VN.n835 VN.n834 0.00946797
R11838 VN.n365 VN.n338 0.00946797
R11839 VN.n297 VN.n296 0.00946797
R11840 VN.n262 VN.n180 0.00946797
R11841 VN.n213 VN.n212 0.00946797
R11842 VN.n416 VN.n393 0.00946797
R11843 VN.n451 VN.n450 0.00946797
R11844 VN.n472 VN.n121 0.00946797
R11845 VN.n86 VN.n74 0.00946797
R11846 VN.n597 VN.n595 0.00946797
R11847 VN.n669 VN.n668 0.00946797
R11848 VN.n699 VN.n554 0.00946797
R11849 VN.n513 VN.n512 0.00946797
R11850 VN.n739 VN.n727 0.00946797
R11851 VN.n813 VN.n793 0.00946797
R11852 VN.n55 VN.n54 0.0088274
R11853 VN.n841 VN.n840 0.0088274
R11854 VN.n373 VN.n333 0.0088274
R11855 VN.n288 VN.n287 0.0088274
R11856 VN.n253 VN.n184 0.0088274
R11857 VN.n203 VN.n202 0.0088274
R11858 VN.n421 VN.n389 0.0088274
R11859 VN.n457 VN.n456 0.0088274
R11860 VN.n478 VN.n477 0.0088274
R11861 VN.n78 VN.n76 0.0088274
R11862 VN.n592 VN.n590 0.0088274
R11863 VN.n678 VN.n677 0.0088274
R11864 VN.n707 VN.n549 0.0088274
R11865 VN.n504 VN.n503 0.0088274
R11866 VN.n730 VN.n729 0.0088274
R11867 VN.n819 VN.n818 0.0088274
R11868 VN.n36 VN.n35 0.00818683
R11869 VN.n786 VN.n784 0.00818683
R11870 VN.n404 VN.n403 0.00818683
R11871 VN.n381 VN.n149 0.00818683
R11872 VN.n133 VN.n131 0.00818683
R11873 VN.n100 VN.n99 0.00818683
R11874 VN.n754 VN.n753 0.00818683
R11875 VN.n804 VN.n0 0.00818683
R11876 VN.n353 VN.n346 0.00690569
R11877 VN.n352 VN.n347 0.00690569
R11878 VN.n312 VN.n311 0.00690569
R11879 VN.n315 VN.n158 0.00690569
R11880 VN.n277 VN.n174 0.00690569
R11881 VN.n279 VN.n278 0.00690569
R11882 VN.n228 VN.n227 0.00690569
R11883 VN.n230 VN.n229 0.00690569
R11884 VN.n605 VN.n603 0.00690569
R11885 VN.n609 VN.n608 0.00690569
R11886 VN.n655 VN.n654 0.00690569
R11887 VN.n651 VN.n579 0.00690569
R11888 VN.n687 VN.n562 0.00690569
R11889 VN.n686 VN.n563 0.00690569
R11890 VN.n528 VN.n527 0.00690569
R11891 VN.n531 VN.n491 0.00690569
R11892 VN VN.n849 0.00306228
R11893 VN.n386 VN.n384 0.00185849
R11894 VN.n428 VN.n387 0.00185849
R11895 VN.n108 VN.n107 0.00185849
R11896 VN.n114 VN.n113 0.00185849
R11897 VN.n13 VN.n12 0.00185849
R11898 VN.n19 VN.n18 0.00185849
R11899 VN.n762 VN.n761 0.00185849
R11900 VN.n768 VN.n767 0.00185849
R11901 VN.n333 VN.n152 0.00178114
R11902 VN.n338 VN.n336 0.00178114
R11903 VN.n343 VN.n341 0.00178114
R11904 VN.n349 VN.n347 0.00178114
R11905 VN.n287 VN.n286 0.00178114
R11906 VN.n296 VN.n295 0.00178114
R11907 VN.n305 VN.n304 0.00178114
R11908 VN.n316 VN.n315 0.00178114
R11909 VN.n249 VN.n184 0.00178114
R11910 VN.n258 VN.n180 0.00178114
R11911 VN.n268 VN.n267 0.00178114
R11912 VN.n278 VN.n172 0.00178114
R11913 VN.n324 VN.n323 0.00178114
R11914 VN.n330 VN.n329 0.00178114
R11915 VN.n240 VN.n239 0.00178114
R11916 VN.n246 VN.n245 0.00178114
R11917 VN.n212 VN.n211 0.00178114
R11918 VN.n219 VN.n194 0.00178114
R11919 VN.n230 VN.n190 0.00178114
R11920 VN.n633 VN.n590 0.00178114
R11921 VN.n625 VN.n595 0.00178114
R11922 VN.n617 VN.n600 0.00178114
R11923 VN.n608 VN.n606 0.00178114
R11924 VN.n679 VN.n678 0.00178114
R11925 VN.n670 VN.n669 0.00178114
R11926 VN.n661 VN.n660 0.00178114
R11927 VN.n651 VN.n650 0.00178114
R11928 VN.n549 VN.n485 0.00178114
R11929 VN.n554 VN.n552 0.00178114
R11930 VN.n559 VN.n557 0.00178114
R11931 VN.n566 VN.n563 0.00178114
R11932 VN.n585 VN.n583 0.00178114
R11933 VN.n638 VN.n586 0.00178114
R11934 VN.n540 VN.n539 0.00178114
R11935 VN.n546 VN.n545 0.00178114
R11936 VN.n512 VN.n511 0.00178114
R11937 VN.n521 VN.n520 0.00178114
R11938 VN.n532 VN.n531 0.00178114
R11939 a_n13990_n5465.n115 a_n13990_n5465.n114 9.23995
R11940 a_n13990_n5465.n24 a_n13990_n5465.n21 7.94229
R11941 a_n13990_n5465.n144 a_n13990_n5465.n142 7.94229
R11942 a_n13990_n5465.n113 a_n13990_n5465.t137 6.72766
R11943 a_n13990_n5465.n95 a_n13990_n5465.n92 6.58329
R11944 a_n13990_n5465.n119 a_n13990_n5465.n115 6.01251
R11945 a_n13990_n5465.n94 a_n13990_n5465.t21 5.85326
R11946 a_n13990_n5465.n90 a_n13990_n5465.t114 5.85326
R11947 a_n13990_n5465.n94 a_n13990_n5465.n93 5.84661
R11948 a_n13990_n5465.n20 a_n13990_n5465.t93 5.69423
R11949 a_n13990_n5465.n25 a_n13990_n5465.t61 5.69423
R11950 a_n13990_n5465.n141 a_n13990_n5465.t62 5.69423
R11951 a_n13990_n5465.n145 a_n13990_n5465.t73 5.69423
R11952 a_n13990_n5465.n20 a_n13990_n5465.n19 5.49558
R11953 a_n13990_n5465.n141 a_n13990_n5465.n140 5.49558
R11954 a_n13990_n5465.n0 a_n13990_n5465.n149 4.22068
R11955 a_n13990_n5465.t30 a_n13990_n5465.n1 5.69068
R11956 a_n13990_n5465.n148 a_n13990_n5465.n2 4.22068
R11957 a_n13990_n5465.n3 a_n13990_n5465.n117 4.22068
R11958 a_n13990_n5465.t48 a_n13990_n5465.n4 5.69068
R11959 a_n13990_n5465.n116 a_n13990_n5465.n5 4.22068
R11960 a_n13990_n5465.n7 a_n13990_n5465.n61 4.58971
R11961 a_n13990_n5465.n8 a_n13990_n5465.t117 5.84971
R11962 a_n13990_n5465.n9 a_n13990_n5465.n66 4.58971
R11963 a_n13990_n5465.n6 a_n13990_n5465.t126 5.47076
R11964 a_n13990_n5465.n92 a_n13990_n5465.n91 4.59326
R11965 a_n13990_n5465.n114 a_n13990_n5465.n113 4.52463
R11966 a_n13990_n5465.n100 a_n13990_n5465.t132 4.41563
R11967 a_n13990_n5465.n109 a_n13990_n5465.t129 4.41563
R11968 a_n13990_n5465.n24 a_n13990_n5465.n23 4.22423
R11969 a_n13990_n5465.n144 a_n13990_n5465.n143 4.22423
R11970 a_n13990_n5465.n113 a_n13990_n5465.n112 4.21432
R11971 a_n13990_n5465.n84 a_n13990_n5465.t5 4.21195
R11972 a_n13990_n5465.n86 a_n13990_n5465.t4 4.21195
R11973 a_n13990_n5465.n71 a_n13990_n5465.t15 4.21195
R11974 a_n13990_n5465.n69 a_n13990_n5465.t0 4.21195
R11975 a_n13990_n5465.n10 a_n13990_n5465.t99 4.05054
R11976 a_n13990_n5465.n154 a_n13990_n5465.t60 4.05054
R11977 a_n13990_n5465.n31 a_n13990_n5465.t41 4.05054
R11978 a_n13990_n5465.n33 a_n13990_n5465.t49 4.05054
R11979 a_n13990_n5465.n39 a_n13990_n5465.t79 4.05054
R11980 a_n13990_n5465.n41 a_n13990_n5465.t92 4.05054
R11981 a_n13990_n5465.n26 a_n13990_n5465.t53 4.05054
R11982 a_n13990_n5465.n51 a_n13990_n5465.t100 4.05054
R11983 a_n13990_n5465.n56 a_n13990_n5465.t111 4.05054
R11984 a_n13990_n5465.n58 a_n13990_n5465.t84 4.05054
R11985 a_n13990_n5465.n126 a_n13990_n5465.t71 4.05054
R11986 a_n13990_n5465.n128 a_n13990_n5465.t45 4.05054
R11987 a_n13990_n5465.n134 a_n13990_n5465.t31 4.05054
R11988 a_n13990_n5465.n136 a_n13990_n5465.t67 4.05054
R11989 a_n13990_n5465.n46 a_n13990_n5465.t36 4.05054
R11990 a_n13990_n5465.t112 a_n13990_n5465.n157 4.05054
R11991 a_n13990_n5465.n84 a_n13990_n5465.t18 4.03668
R11992 a_n13990_n5465.n86 a_n13990_n5465.t23 4.03668
R11993 a_n13990_n5465.n71 a_n13990_n5465.t8 4.03668
R11994 a_n13990_n5465.n69 a_n13990_n5465.t11 4.03668
R11995 a_n13990_n5465.n157 a_n13990_n5465.t110 3.87765
R11996 a_n13990_n5465.n10 a_n13990_n5465.t98 3.87765
R11997 a_n13990_n5465.n154 a_n13990_n5465.t58 3.87765
R11998 a_n13990_n5465.n31 a_n13990_n5465.t40 3.87765
R11999 a_n13990_n5465.n33 a_n13990_n5465.t46 3.87765
R12000 a_n13990_n5465.n39 a_n13990_n5465.t78 3.87765
R12001 a_n13990_n5465.n41 a_n13990_n5465.t91 3.87765
R12002 a_n13990_n5465.n26 a_n13990_n5465.t52 3.87765
R12003 a_n13990_n5465.n51 a_n13990_n5465.t103 3.87765
R12004 a_n13990_n5465.n56 a_n13990_n5465.t25 3.87765
R12005 a_n13990_n5465.n58 a_n13990_n5465.t86 3.87765
R12006 a_n13990_n5465.n126 a_n13990_n5465.t72 3.87765
R12007 a_n13990_n5465.n128 a_n13990_n5465.t47 3.87765
R12008 a_n13990_n5465.n134 a_n13990_n5465.t33 3.87765
R12009 a_n13990_n5465.n136 a_n13990_n5465.t68 3.87765
R12010 a_n13990_n5465.n46 a_n13990_n5465.t38 3.87765
R12011 a_n13990_n5465.n100 a_n13990_n5465.t133 3.833
R12012 a_n13990_n5465.n109 a_n13990_n5465.t128 3.833
R12013 a_n13990_n5465.n80 a_n13990_n5465.n76 3.81703
R12014 a_n13990_n5465.n67 a_n13990_n5465.n9 3.95161
R12015 a_n13990_n5465.n108 a_n13990_n5465.n104 3.80578
R12016 a_n13990_n5465.n99 a_n13990_n5465.n6 3.90344
R12017 a_n13990_n5465.n97 a_n13990_n5465.n96 3.69568
R12018 a_n13990_n5465.n44 a_n13990_n5465.n25 3.25667
R12019 a_n13990_n5465.n103 a_n13990_n5465.n101 3.15563
R12020 a_n13990_n5465.n107 a_n13990_n5465.n105 3.15563
R12021 a_n13990_n5465.n2 a_n13990_n5465.n147 3.15553
R12022 a_n13990_n5465.n5 a_n13990_n5465.n45 3.15553
R12023 a_n13990_n5465.n83 a_n13990_n5465.n82 2.95195
R12024 a_n13990_n5465.n79 a_n13990_n5465.n78 2.95195
R12025 a_n13990_n5465.n75 a_n13990_n5465.n74 2.95195
R12026 a_n13990_n5465.n65 a_n13990_n5465.n64 2.95195
R12027 a_n13990_n5465.n83 a_n13990_n5465.n81 2.77668
R12028 a_n13990_n5465.n79 a_n13990_n5465.n77 2.77668
R12029 a_n13990_n5465.n75 a_n13990_n5465.n73 2.77668
R12030 a_n13990_n5465.n65 a_n13990_n5465.n63 2.77668
R12031 a_n13990_n5465.n50 a_n13990_n5465.n46 2.73714
R12032 a_n13990_n5465.n30 a_n13990_n5465.n26 2.73714
R12033 a_n13990_n5465.n14 a_n13990_n5465.n10 2.73672
R12034 a_n13990_n5465.n55 a_n13990_n5465.n51 2.73672
R12035 a_n13990_n5465.n104 a_n13990_n5465.n100 2.71872
R12036 a_n13990_n5465.n85 a_n13990_n5465.n83 2.71872
R12037 a_n13990_n5465.n129 a_n13990_n5465.n127 2.60203
R12038 a_n13990_n5465.n34 a_n13990_n5465.n32 2.60203
R12039 a_n13990_n5465.n97 a_n13990_n5465.n60 2.5825
R12040 a_n13990_n5465.n13 a_n13990_n5465.n12 2.58054
R12041 a_n13990_n5465.n17 a_n13990_n5465.n16 2.58054
R12042 a_n13990_n5465.n37 a_n13990_n5465.n36 2.58054
R12043 a_n13990_n5465.n29 a_n13990_n5465.n28 2.58054
R12044 a_n13990_n5465.n54 a_n13990_n5465.n53 2.58054
R12045 a_n13990_n5465.n124 a_n13990_n5465.n123 2.58054
R12046 a_n13990_n5465.n132 a_n13990_n5465.n131 2.58054
R12047 a_n13990_n5465.n49 a_n13990_n5465.n48 2.58054
R12048 a_n13990_n5465.n103 a_n13990_n5465.n102 2.573
R12049 a_n13990_n5465.n107 a_n13990_n5465.n106 2.573
R12050 a_n13990_n5465.n72 a_n13990_n5465.n70 2.56118
R12051 a_n13990_n5465.n87 a_n13990_n5465.n85 2.56118
R12052 a_n13990_n5465.n90 a_n13990_n5465.n60 2.54573
R12053 a_n13990_n5465.n137 a_n13990_n5465.n135 2.53418
R12054 a_n13990_n5465.n59 a_n13990_n5465.n57 2.53418
R12055 a_n13990_n5465.n42 a_n13990_n5465.n40 2.53418
R12056 a_n13990_n5465.n156 a_n13990_n5465.n155 2.53418
R12057 a_n13990_n5465.n146 a_n13990_n5465.n145 2.51873
R12058 a_n13990_n5465.n13 a_n13990_n5465.n11 2.40765
R12059 a_n13990_n5465.n17 a_n13990_n5465.n15 2.40765
R12060 a_n13990_n5465.n37 a_n13990_n5465.n35 2.40765
R12061 a_n13990_n5465.n29 a_n13990_n5465.n27 2.40765
R12062 a_n13990_n5465.n54 a_n13990_n5465.n52 2.40765
R12063 a_n13990_n5465.n124 a_n13990_n5465.n122 2.40765
R12064 a_n13990_n5465.n132 a_n13990_n5465.n130 2.40765
R12065 a_n13990_n5465.n49 a_n13990_n5465.n47 2.40765
R12066 a_n13990_n5465.n89 a_n13990_n5465.n62 2.27857
R12067 a_n13990_n5465.n152 a_n13990_n5465.n21 2.23844
R12068 a_n13990_n5465.n68 a_n13990_n5465.n65 2.00466
R12069 a_n13990_n5465.n111 a_n13990_n5465.n110 1.67718
R12070 a_n13990_n5465.n62 a_n13990_n5465.n7 1.67353
R12071 a_n13990_n5465.n150 a_n13990_n5465.n0 1.65553
R12072 a_n13990_n5465.n118 a_n13990_n5465.n3 1.65553
R12073 a_n13990_n5465.n139 a_n13990_n5465.n138 1.5005
R12074 a_n13990_n5465.n68 a_n13990_n5465.n67 1.5005
R12075 a_n13990_n5465.n89 a_n13990_n5465.n88 1.5005
R12076 a_n13990_n5465.n96 a_n13990_n5465.n95 1.5005
R12077 a_n13990_n5465.n119 a_n13990_n5465.n118 1.5005
R12078 a_n13990_n5465.n121 a_n13990_n5465.n120 1.5005
R12079 a_n13990_n5465.n142 a_n13990_n5465.n22 1.5005
R12080 a_n13990_n5465.n151 a_n13990_n5465.n150 1.5005
R12081 a_n13990_n5465.n153 a_n13990_n5465.n152 1.5005
R12082 a_n13990_n5465.n44 a_n13990_n5465.n43 1.5005
R12083 a_n13990_n5465.n11 a_n13990_n5465.t27 1.4705
R12084 a_n13990_n5465.n11 a_n13990_n5465.t74 1.4705
R12085 a_n13990_n5465.n12 a_n13990_n5465.t29 1.4705
R12086 a_n13990_n5465.n12 a_n13990_n5465.t75 1.4705
R12087 a_n13990_n5465.n15 a_n13990_n5465.t101 1.4705
R12088 a_n13990_n5465.n15 a_n13990_n5465.t81 1.4705
R12089 a_n13990_n5465.n16 a_n13990_n5465.t105 1.4705
R12090 a_n13990_n5465.n16 a_n13990_n5465.t82 1.4705
R12091 a_n13990_n5465.n35 a_n13990_n5465.t83 1.4705
R12092 a_n13990_n5465.n35 a_n13990_n5465.t37 1.4705
R12093 a_n13990_n5465.n36 a_n13990_n5465.t85 1.4705
R12094 a_n13990_n5465.n36 a_n13990_n5465.t39 1.4705
R12095 a_n13990_n5465.n27 a_n13990_n5465.t42 1.4705
R12096 a_n13990_n5465.n27 a_n13990_n5465.t34 1.4705
R12097 a_n13990_n5465.n28 a_n13990_n5465.t44 1.4705
R12098 a_n13990_n5465.n28 a_n13990_n5465.t35 1.4705
R12099 a_n13990_n5465.n19 a_n13990_n5465.t32 1.4705
R12100 a_n13990_n5465.n19 a_n13990_n5465.t94 1.4705
R12101 a_n13990_n5465.n23 a_n13990_n5465.t70 1.4705
R12102 a_n13990_n5465.n23 a_n13990_n5465.t43 1.4705
R12103 a_n13990_n5465.n149 a_n13990_n5465.t69 1.4705
R12104 a_n13990_n5465.n149 a_n13990_n5465.t95 1.4705
R12105 a_n13990_n5465.n148 a_n13990_n5465.t28 1.4705
R12106 a_n13990_n5465.n148 a_n13990_n5465.t66 1.4705
R12107 a_n13990_n5465.n140 a_n13990_n5465.t59 1.4705
R12108 a_n13990_n5465.n140 a_n13990_n5465.t88 1.4705
R12109 a_n13990_n5465.n143 a_n13990_n5465.t87 1.4705
R12110 a_n13990_n5465.n143 a_n13990_n5465.t26 1.4705
R12111 a_n13990_n5465.n52 a_n13990_n5465.t51 1.4705
R12112 a_n13990_n5465.n52 a_n13990_n5465.t107 1.4705
R12113 a_n13990_n5465.n53 a_n13990_n5465.t50 1.4705
R12114 a_n13990_n5465.n53 a_n13990_n5465.t106 1.4705
R12115 a_n13990_n5465.n122 a_n13990_n5465.t97 1.4705
R12116 a_n13990_n5465.n122 a_n13990_n5465.t57 1.4705
R12117 a_n13990_n5465.n123 a_n13990_n5465.t96 1.4705
R12118 a_n13990_n5465.n123 a_n13990_n5465.t56 1.4705
R12119 a_n13990_n5465.n130 a_n13990_n5465.t55 1.4705
R12120 a_n13990_n5465.n130 a_n13990_n5465.t109 1.4705
R12121 a_n13990_n5465.n131 a_n13990_n5465.t54 1.4705
R12122 a_n13990_n5465.n131 a_n13990_n5465.t108 1.4705
R12123 a_n13990_n5465.n47 a_n13990_n5465.t90 1.4705
R12124 a_n13990_n5465.n47 a_n13990_n5465.t65 1.4705
R12125 a_n13990_n5465.n48 a_n13990_n5465.t89 1.4705
R12126 a_n13990_n5465.n48 a_n13990_n5465.t63 1.4705
R12127 a_n13990_n5465.n117 a_n13990_n5465.t77 1.4705
R12128 a_n13990_n5465.n117 a_n13990_n5465.t76 1.4705
R12129 a_n13990_n5465.n116 a_n13990_n5465.t80 1.4705
R12130 a_n13990_n5465.n116 a_n13990_n5465.t102 1.4705
R12131 a_n13990_n5465.n14 a_n13990_n5465.n13 1.46537
R12132 a_n13990_n5465.n157 a_n13990_n5465.n156 1.46537
R12133 a_n13990_n5465.n18 a_n13990_n5465.n17 1.46537
R12134 a_n13990_n5465.n32 a_n13990_n5465.n31 1.46537
R12135 a_n13990_n5465.n34 a_n13990_n5465.n33 1.46537
R12136 a_n13990_n5465.n38 a_n13990_n5465.n37 1.46537
R12137 a_n13990_n5465.n40 a_n13990_n5465.n39 1.46537
R12138 a_n13990_n5465.n30 a_n13990_n5465.n29 1.46537
R12139 a_n13990_n5465.n55 a_n13990_n5465.n54 1.46537
R12140 a_n13990_n5465.n57 a_n13990_n5465.n56 1.46537
R12141 a_n13990_n5465.n125 a_n13990_n5465.n124 1.46537
R12142 a_n13990_n5465.n127 a_n13990_n5465.n126 1.46537
R12143 a_n13990_n5465.n129 a_n13990_n5465.n128 1.46537
R12144 a_n13990_n5465.n133 a_n13990_n5465.n132 1.46537
R12145 a_n13990_n5465.n135 a_n13990_n5465.n134 1.46537
R12146 a_n13990_n5465.n50 a_n13990_n5465.n49 1.46537
R12147 a_n13990_n5465.n85 a_n13990_n5465.n84 1.46537
R12148 a_n13990_n5465.n80 a_n13990_n5465.n79 1.46537
R12149 a_n13990_n5465.n76 a_n13990_n5465.n75 1.46537
R12150 a_n13990_n5465.n72 a_n13990_n5465.n71 1.46537
R12151 a_n13990_n5465.n104 a_n13990_n5465.n103 1.46537
R12152 a_n13990_n5465.n108 a_n13990_n5465.n107 1.46537
R12153 a_n13990_n5465.n110 a_n13990_n5465.n109 1.46537
R12154 a_n13990_n5465.n155 a_n13990_n5465.n154 1.46535
R12155 a_n13990_n5465.n42 a_n13990_n5465.n41 1.46535
R12156 a_n13990_n5465.n59 a_n13990_n5465.n58 1.46535
R12157 a_n13990_n5465.n137 a_n13990_n5465.n136 1.46535
R12158 a_n13990_n5465.n87 a_n13990_n5465.n86 1.46535
R12159 a_n13990_n5465.n70 a_n13990_n5465.n69 1.46535
R12160 a_n13990_n5465.n115 a_n13990_n5465.n45 1.43535
R12161 a_n13990_n5465.n99 a_n13990_n5465.n97 1.31908
R12162 a_n13990_n5465.n156 a_n13990_n5465.n14 1.27228
R12163 a_n13990_n5465.n25 a_n13990_n5465.n24 1.27228
R12164 a_n13990_n5465.n145 a_n13990_n5465.n144 1.27228
R12165 a_n13990_n5465.n135 a_n13990_n5465.n133 1.27228
R12166 a_n13990_n5465.n133 a_n13990_n5465.n129 1.27228
R12167 a_n13990_n5465.n127 a_n13990_n5465.n125 1.27228
R12168 a_n13990_n5465.n57 a_n13990_n5465.n55 1.27228
R12169 a_n13990_n5465.n40 a_n13990_n5465.n38 1.27228
R12170 a_n13990_n5465.n38 a_n13990_n5465.n34 1.27228
R12171 a_n13990_n5465.n32 a_n13990_n5465.n18 1.27228
R12172 a_n13990_n5465.n101 a_n13990_n5465.t121 1.2605
R12173 a_n13990_n5465.n101 a_n13990_n5465.t130 1.2605
R12174 a_n13990_n5465.n102 a_n13990_n5465.t134 1.2605
R12175 a_n13990_n5465.n102 a_n13990_n5465.t131 1.2605
R12176 a_n13990_n5465.n105 a_n13990_n5465.t123 1.2605
R12177 a_n13990_n5465.n105 a_n13990_n5465.t136 1.2605
R12178 a_n13990_n5465.n106 a_n13990_n5465.t135 1.2605
R12179 a_n13990_n5465.n106 a_n13990_n5465.t127 1.2605
R12180 a_n13990_n5465.n112 a_n13990_n5465.t138 1.2605
R12181 a_n13990_n5465.n112 a_n13990_n5465.t122 1.2605
R12182 a_n13990_n5465.n98 a_n13990_n5465.t124 1.2605
R12183 a_n13990_n5465.n98 a_n13990_n5465.t125 1.2605
R12184 a_n13990_n5465.n61 a_n13990_n5465.t119 1.2605
R12185 a_n13990_n5465.n61 a_n13990_n5465.t17 1.2605
R12186 a_n13990_n5465.n66 a_n13990_n5465.t116 1.2605
R12187 a_n13990_n5465.n66 a_n13990_n5465.t140 1.2605
R12188 a_n13990_n5465.n93 a_n13990_n5465.t14 1.2605
R12189 a_n13990_n5465.n93 a_n13990_n5465.t10 1.2605
R12190 a_n13990_n5465.n91 a_n13990_n5465.t2 1.2605
R12191 a_n13990_n5465.n91 a_n13990_n5465.t115 1.2605
R12192 a_n13990_n5465.n81 a_n13990_n5465.t13 1.2605
R12193 a_n13990_n5465.n81 a_n13990_n5465.t19 1.2605
R12194 a_n13990_n5465.n82 a_n13990_n5465.t20 1.2605
R12195 a_n13990_n5465.n82 a_n13990_n5465.t6 1.2605
R12196 a_n13990_n5465.n77 a_n13990_n5465.t113 1.2605
R12197 a_n13990_n5465.n77 a_n13990_n5465.t7 1.2605
R12198 a_n13990_n5465.n78 a_n13990_n5465.t118 1.2605
R12199 a_n13990_n5465.n78 a_n13990_n5465.t24 1.2605
R12200 a_n13990_n5465.n73 a_n13990_n5465.t3 1.2605
R12201 a_n13990_n5465.n73 a_n13990_n5465.t9 1.2605
R12202 a_n13990_n5465.n74 a_n13990_n5465.t1 1.2605
R12203 a_n13990_n5465.n74 a_n13990_n5465.t16 1.2605
R12204 a_n13990_n5465.n63 a_n13990_n5465.t141 1.2605
R12205 a_n13990_n5465.n63 a_n13990_n5465.t22 1.2605
R12206 a_n13990_n5465.n64 a_n13990_n5465.t139 1.2605
R12207 a_n13990_n5465.n64 a_n13990_n5465.t12 1.2605
R12208 a_n13990_n5465.n92 a_n13990_n5465.n90 1.25428
R12209 a_n13990_n5465.n76 a_n13990_n5465.n72 1.25428
R12210 a_n13990_n5465.n110 a_n13990_n5465.n108 1.25428
R12211 a_n13990_n5465.n95 a_n13990_n5465.n94 1.04573
R12212 a_n13990_n5465.n21 a_n13990_n5465.n20 1.01873
R12213 a_n13990_n5465.n142 a_n13990_n5465.n141 1.01873
R12214 a_n13990_n5465.n147 a_n13990_n5465.n44 0.778574
R12215 a_n13990_n5465.n139 a_n13990_n5465.n45 0.778574
R12216 a_n13990_n5465.n152 a_n13990_n5465.n151 0.778574
R12217 a_n13990_n5465.n120 a_n13990_n5465.n119 0.778574
R12218 a_n13990_n5465.n146 a_n13990_n5465.n139 0.738439
R12219 a_n13990_n5465.n67 a_n13990_n5465.n60 0.738439
R12220 a_n13990_n5465.n96 a_n13990_n5465.n89 0.738439
R12221 a_n13990_n5465.n120 a_n13990_n5465.n22 0.738439
R12222 a_n13990_n5465.n114 a_n13990_n5465.n111 0.737223
R12223 a_n13990_n5465.n138 a_n13990_n5465.n137 0.699581
R12224 a_n13990_n5465.n121 a_n13990_n5465.n59 0.699581
R12225 a_n13990_n5465.n70 a_n13990_n5465.n68 0.699581
R12226 a_n13990_n5465.n88 a_n13990_n5465.n87 0.699581
R12227 a_n13990_n5465.n43 a_n13990_n5465.n42 0.699581
R12228 a_n13990_n5465.n155 a_n13990_n5465.n153 0.699581
R12229 a_n13990_n5465.n111 a_n13990_n5465.n99 0.585196
R12230 a_n13990_n5465.n138 a_n13990_n5465.n50 0.557791
R12231 a_n13990_n5465.n125 a_n13990_n5465.n121 0.557791
R12232 a_n13990_n5465.n43 a_n13990_n5465.n30 0.557791
R12233 a_n13990_n5465.n153 a_n13990_n5465.n18 0.557791
R12234 a_n13990_n5465.n88 a_n13990_n5465.n80 0.539791
R12235 a_n13990_n5465.n147 a_n13990_n5465.n146 0.530466
R12236 a_n13990_n5465.n151 a_n13990_n5465.n22 0.530466
R12237 a_n13990_n5465.n1 a_n13990_n5465.n2 1.27228
R12238 a_n13990_n5465.n150 a_n13990_n5465.n1 7.30549
R12239 a_n13990_n5465.t64 a_n13990_n5465.n0 6.96214
R12240 a_n13990_n5465.n4 a_n13990_n5465.n5 1.27228
R12241 a_n13990_n5465.n118 a_n13990_n5465.n4 7.30549
R12242 a_n13990_n5465.t104 a_n13990_n5465.n3 6.96214
R12243 a_n13990_n5465.n98 a_n13990_n5465.n6 5.45652
R12244 a_n13990_n5465.n8 a_n13990_n5465.n9 1.25428
R12245 a_n13990_n5465.n62 a_n13990_n5465.n8 5.95549
R12246 a_n13990_n5465.t120 a_n13990_n5465.n7 7.10317
R12247 a_5396_9163.n33 a_5396_9163.n30 7.94229
R12248 a_5396_9163.n74 a_5396_9163.n72 7.94229
R12249 a_5396_9163.n98 a_5396_9163.t168 6.58663
R12250 a_5396_9163.n138 a_5396_9163.t109 6.58663
R12251 a_5396_9163.n184 a_5396_9163.n183 5.95439
R12252 a_5396_9163.n140 a_5396_9163.n139 5.95439
R12253 a_5396_9163.n32 a_5396_9163.t19 5.69423
R12254 a_5396_9163.n28 a_5396_9163.t33 5.69423
R12255 a_5396_9163.n71 a_5396_9163.t57 5.69423
R12256 a_5396_9163.n75 a_5396_9163.t67 5.69423
R12257 a_5396_9163.n32 a_5396_9163.n31 5.49558
R12258 a_5396_9163.n71 a_5396_9163.n70 5.49558
R12259 a_5396_9163.n184 a_5396_9163.t118 5.31528
R12260 a_5396_9163.n140 a_5396_9163.t112 5.31528
R12261 a_5396_9163.n0 a_5396_9163.n27 4.22068
R12262 a_5396_9163.n1 a_5396_9163.t82 5.69068
R12263 a_5396_9163.n2 a_5396_9163.n26 4.22068
R12264 a_5396_9163.n3 a_5396_9163.n191 4.22068
R12265 a_5396_9163.t13 a_5396_9163.n4 5.69068
R12266 a_5396_9163.n190 a_5396_9163.n5 4.22068
R12267 a_5396_9163.n115 a_5396_9163.n7 3.84173
R12268 a_5396_9163.n145 a_5396_9163.n10 3.84173
R12269 a_5396_9163.n6 a_5396_9163.t120 5.31173
R12270 a_5396_9163.t145 a_5396_9163.n8 5.31173
R12271 a_5396_9163.n9 a_5396_9163.t173 5.31173
R12272 a_5396_9163.t104 a_5396_9163.n11 5.31173
R12273 a_5396_9163.n187 a_5396_9163.n186 4.50663
R12274 a_5396_9163.n143 a_5396_9163.n142 4.50663
R12275 a_5396_9163.n136 a_5396_9163.n8 4.46113
R12276 a_5396_9163.n30 a_5396_9163.n29 4.22423
R12277 a_5396_9163.n74 a_5396_9163.n73 4.22423
R12278 a_5396_9163.n12 a_5396_9163.t84 4.05054
R12279 a_5396_9163.n17 a_5396_9163.t14 4.05054
R12280 a_5396_9163.n82 a_5396_9163.t70 4.05054
R12281 a_5396_9163.n84 a_5396_9163.t46 4.05054
R12282 a_5396_9163.n90 a_5396_9163.t85 4.05054
R12283 a_5396_9163.n92 a_5396_9163.t52 4.05054
R12284 a_5396_9163.n77 a_5396_9163.t24 4.05054
R12285 a_5396_9163.n56 a_5396_9163.t42 4.05054
R12286 a_5396_9163.n61 a_5396_9163.t61 4.05054
R12287 a_5396_9163.n63 a_5396_9163.t18 4.05054
R12288 a_5396_9163.n50 a_5396_9163.t5 4.05054
R12289 a_5396_9163.n48 a_5396_9163.t54 4.05054
R12290 a_5396_9163.n42 a_5396_9163.t51 4.05054
R12291 a_5396_9163.n40 a_5396_9163.t28 4.05054
R12292 a_5396_9163.n34 a_5396_9163.t86 4.05054
R12293 a_5396_9163.t87 a_5396_9163.n197 4.05054
R12294 a_5396_9163.n188 a_5396_9163.n24 3.97558
R12295 a_5396_9163.n197 a_5396_9163.t50 3.87765
R12296 a_5396_9163.n12 a_5396_9163.t73 3.87765
R12297 a_5396_9163.n17 a_5396_9163.t4 3.87765
R12298 a_5396_9163.n82 a_5396_9163.t37 3.87765
R12299 a_5396_9163.n84 a_5396_9163.t83 3.87765
R12300 a_5396_9163.n90 a_5396_9163.t79 3.87765
R12301 a_5396_9163.n92 a_5396_9163.t59 3.87765
R12302 a_5396_9163.n77 a_5396_9163.t30 3.87765
R12303 a_5396_9163.n56 a_5396_9163.t35 3.87765
R12304 a_5396_9163.n61 a_5396_9163.t55 3.87765
R12305 a_5396_9163.n63 a_5396_9163.t10 3.87765
R12306 a_5396_9163.n50 a_5396_9163.t0 3.87765
R12307 a_5396_9163.n48 a_5396_9163.t49 3.87765
R12308 a_5396_9163.n42 a_5396_9163.t47 3.87765
R12309 a_5396_9163.n40 a_5396_9163.t22 3.87765
R12310 a_5396_9163.n34 a_5396_9163.t78 3.87765
R12311 a_5396_9163.n98 a_5396_9163.n97 3.84528
R12312 a_5396_9163.n186 a_5396_9163.n185 3.84528
R12313 a_5396_9163.n138 a_5396_9163.n137 3.84528
R12314 a_5396_9163.n142 a_5396_9163.n141 3.84528
R12315 a_5396_9163.n160 a_5396_9163.n156 3.79678
R12316 a_5396_9163.n175 a_5396_9163.n171 3.79678
R12317 a_5396_9163.n131 a_5396_9163.n127 3.79678
R12318 a_5396_9163.n110 a_5396_9163.n106 3.79678
R12319 a_5396_9163.n11 a_5396_9163.n144 3.87644
R12320 a_5396_9163.n180 a_5396_9163.n164 3.73034
R12321 a_5396_9163.n123 a_5396_9163.n119 3.73034
R12322 a_5396_9163.n28 a_5396_9163.n25 3.25667
R12323 a_5396_9163.n69 a_5396_9163.n2 3.15553
R12324 a_5396_9163.n5 a_5396_9163.n189 3.15553
R12325 a_5396_9163.n183 a_5396_9163.n98 3.00663
R12326 a_5396_9163.n139 a_5396_9163.n138 3.00663
R12327 a_5396_9163.n167 a_5396_9163.n165 2.7866
R12328 a_5396_9163.n170 a_5396_9163.n168 2.7866
R12329 a_5396_9163.n174 a_5396_9163.n172 2.7866
R12330 a_5396_9163.n178 a_5396_9163.n176 2.7866
R12331 a_5396_9163.n163 a_5396_9163.n161 2.7866
R12332 a_5396_9163.n159 a_5396_9163.n157 2.7866
R12333 a_5396_9163.n155 a_5396_9163.n153 2.7866
R12334 a_5396_9163.n151 a_5396_9163.n149 2.7866
R12335 a_5396_9163.n102 a_5396_9163.n100 2.7866
R12336 a_5396_9163.n105 a_5396_9163.n103 2.7866
R12337 a_5396_9163.n109 a_5396_9163.n107 2.7866
R12338 a_5396_9163.n113 a_5396_9163.n111 2.7866
R12339 a_5396_9163.n122 a_5396_9163.n120 2.7866
R12340 a_5396_9163.n126 a_5396_9163.n124 2.7866
R12341 a_5396_9163.n130 a_5396_9163.n128 2.7866
R12342 a_5396_9163.n134 a_5396_9163.n132 2.7866
R12343 a_5396_9163.n38 a_5396_9163.n34 2.73714
R12344 a_5396_9163.n81 a_5396_9163.n77 2.73714
R12345 a_5396_9163.n16 a_5396_9163.n12 2.73672
R12346 a_5396_9163.n60 a_5396_9163.n56 2.73672
R12347 a_5396_9163.n171 a_5396_9163.n167 2.73672
R12348 a_5396_9163.n106 a_5396_9163.n102 2.73672
R12349 a_5396_9163.n51 a_5396_9163.n49 2.60203
R12350 a_5396_9163.n85 a_5396_9163.n83 2.60203
R12351 a_5396_9163.n15 a_5396_9163.n14 2.58054
R12352 a_5396_9163.n21 a_5396_9163.n20 2.58054
R12353 a_5396_9163.n88 a_5396_9163.n87 2.58054
R12354 a_5396_9163.n80 a_5396_9163.n79 2.58054
R12355 a_5396_9163.n59 a_5396_9163.n58 2.58054
R12356 a_5396_9163.n54 a_5396_9163.n53 2.58054
R12357 a_5396_9163.n46 a_5396_9163.n45 2.58054
R12358 a_5396_9163.n37 a_5396_9163.n36 2.58054
R12359 a_5396_9163.n196 a_5396_9163.n18 2.53418
R12360 a_5396_9163.n43 a_5396_9163.n41 2.53418
R12361 a_5396_9163.n64 a_5396_9163.n62 2.53418
R12362 a_5396_9163.n93 a_5396_9163.n91 2.53418
R12363 a_5396_9163.n76 a_5396_9163.n75 2.51873
R12364 a_5396_9163.n15 a_5396_9163.n13 2.40765
R12365 a_5396_9163.n21 a_5396_9163.n19 2.40765
R12366 a_5396_9163.n88 a_5396_9163.n86 2.40765
R12367 a_5396_9163.n80 a_5396_9163.n78 2.40765
R12368 a_5396_9163.n59 a_5396_9163.n57 2.40765
R12369 a_5396_9163.n54 a_5396_9163.n52 2.40765
R12370 a_5396_9163.n46 a_5396_9163.n44 2.40765
R12371 a_5396_9163.n37 a_5396_9163.n35 2.40765
R12372 a_5396_9163.n147 a_5396_9163.n9 2.37644
R12373 a_5396_9163.n117 a_5396_9163.n6 2.37644
R12374 a_5396_9163.n66 a_5396_9163.n33 2.23844
R12375 a_5396_9163.n167 a_5396_9163.n166 2.2016
R12376 a_5396_9163.n170 a_5396_9163.n169 2.2016
R12377 a_5396_9163.n174 a_5396_9163.n173 2.2016
R12378 a_5396_9163.n178 a_5396_9163.n177 2.2016
R12379 a_5396_9163.n163 a_5396_9163.n162 2.2016
R12380 a_5396_9163.n159 a_5396_9163.n158 2.2016
R12381 a_5396_9163.n155 a_5396_9163.n154 2.2016
R12382 a_5396_9163.n151 a_5396_9163.n150 2.2016
R12383 a_5396_9163.n102 a_5396_9163.n101 2.2016
R12384 a_5396_9163.n105 a_5396_9163.n104 2.2016
R12385 a_5396_9163.n109 a_5396_9163.n108 2.2016
R12386 a_5396_9163.n113 a_5396_9163.n112 2.2016
R12387 a_5396_9163.n122 a_5396_9163.n121 2.2016
R12388 a_5396_9163.n126 a_5396_9163.n125 2.2016
R12389 a_5396_9163.n130 a_5396_9163.n129 2.2016
R12390 a_5396_9163.n134 a_5396_9163.n133 2.2016
R12391 a_5396_9163.n118 a_5396_9163.n117 2.0852
R12392 a_5396_9163.n188 a_5396_9163.n187 1.85726
R12393 a_5396_9163.n193 a_5396_9163.n24 1.83738
R12394 a_5396_9163.n152 a_5396_9163.n96 1.65018
R12395 a_5396_9163.n136 a_5396_9163.n135 1.65018
R12396 a_5396_9163.n68 a_5396_9163.n0 1.65553
R12397 a_5396_9163.n192 a_5396_9163.n3 1.65553
R12398 a_5396_9163.n39 a_5396_9163.n25 1.5005
R12399 a_5396_9163.n139 a_5396_9163.n99 1.5005
R12400 a_5396_9163.n148 a_5396_9163.n147 1.5005
R12401 a_5396_9163.n183 a_5396_9163.n182 1.5005
R12402 a_5396_9163.n119 a_5396_9163.n118 1.5005
R12403 a_5396_9163.n181 a_5396_9163.n180 1.5005
R12404 a_5396_9163.n193 a_5396_9163.n192 1.5005
R12405 a_5396_9163.n72 a_5396_9163.n23 1.5005
R12406 a_5396_9163.n68 a_5396_9163.n67 1.5005
R12407 a_5396_9163.n66 a_5396_9163.n65 1.5005
R12408 a_5396_9163.n195 a_5396_9163.n194 1.5005
R12409 a_5396_9163.n95 a_5396_9163.n94 1.5005
R12410 a_5396_9163.n13 a_5396_9163.t64 1.4705
R12411 a_5396_9163.n13 a_5396_9163.t44 1.4705
R12412 a_5396_9163.n14 a_5396_9163.t43 1.4705
R12413 a_5396_9163.n14 a_5396_9163.t39 1.4705
R12414 a_5396_9163.n19 a_5396_9163.t16 1.4705
R12415 a_5396_9163.n19 a_5396_9163.t68 1.4705
R12416 a_5396_9163.n20 a_5396_9163.t65 1.4705
R12417 a_5396_9163.n20 a_5396_9163.t2 1.4705
R12418 a_5396_9163.n86 a_5396_9163.t53 1.4705
R12419 a_5396_9163.n86 a_5396_9163.t27 1.4705
R12420 a_5396_9163.n87 a_5396_9163.t25 1.4705
R12421 a_5396_9163.n87 a_5396_9163.t17 1.4705
R12422 a_5396_9163.n78 a_5396_9163.t8 1.4705
R12423 a_5396_9163.n78 a_5396_9163.t75 1.4705
R12424 a_5396_9163.n79 a_5396_9163.t15 1.4705
R12425 a_5396_9163.n79 a_5396_9163.t56 1.4705
R12426 a_5396_9163.n31 a_5396_9163.t77 1.4705
R12427 a_5396_9163.n31 a_5396_9163.t60 1.4705
R12428 a_5396_9163.n29 a_5396_9163.t3 1.4705
R12429 a_5396_9163.n29 a_5396_9163.t72 1.4705
R12430 a_5396_9163.n57 a_5396_9163.t26 1.4705
R12431 a_5396_9163.n57 a_5396_9163.t6 1.4705
R12432 a_5396_9163.n58 a_5396_9163.t32 1.4705
R12433 a_5396_9163.n58 a_5396_9163.t9 1.4705
R12434 a_5396_9163.n52 a_5396_9163.t69 1.4705
R12435 a_5396_9163.n52 a_5396_9163.t34 1.4705
R12436 a_5396_9163.n53 a_5396_9163.t74 1.4705
R12437 a_5396_9163.n53 a_5396_9163.t38 1.4705
R12438 a_5396_9163.n44 a_5396_9163.t12 1.4705
R12439 a_5396_9163.n44 a_5396_9163.t76 1.4705
R12440 a_5396_9163.n45 a_5396_9163.t23 1.4705
R12441 a_5396_9163.n45 a_5396_9163.t80 1.4705
R12442 a_5396_9163.n35 a_5396_9163.t62 1.4705
R12443 a_5396_9163.n35 a_5396_9163.t41 1.4705
R12444 a_5396_9163.n36 a_5396_9163.t66 1.4705
R12445 a_5396_9163.n36 a_5396_9163.t48 1.4705
R12446 a_5396_9163.n27 a_5396_9163.t31 1.4705
R12447 a_5396_9163.n27 a_5396_9163.t1 1.4705
R12448 a_5396_9163.n26 a_5396_9163.t45 1.4705
R12449 a_5396_9163.n26 a_5396_9163.t11 1.4705
R12450 a_5396_9163.n70 a_5396_9163.t29 1.4705
R12451 a_5396_9163.n70 a_5396_9163.t7 1.4705
R12452 a_5396_9163.n73 a_5396_9163.t40 1.4705
R12453 a_5396_9163.n73 a_5396_9163.t20 1.4705
R12454 a_5396_9163.n191 a_5396_9163.t36 1.4705
R12455 a_5396_9163.n191 a_5396_9163.t63 1.4705
R12456 a_5396_9163.n190 a_5396_9163.t81 1.4705
R12457 a_5396_9163.n190 a_5396_9163.t21 1.4705
R12458 a_5396_9163.n116 a_5396_9163.t115 1.4705
R12459 a_5396_9163.n116 a_5396_9163.t113 1.4705
R12460 a_5396_9163.n115 a_5396_9163.t136 1.4705
R12461 a_5396_9163.n115 a_5396_9163.t102 1.4705
R12462 a_5396_9163.n165 a_5396_9163.t94 1.4705
R12463 a_5396_9163.n165 a_5396_9163.t161 1.4705
R12464 a_5396_9163.n166 a_5396_9163.t95 1.4705
R12465 a_5396_9163.n166 a_5396_9163.t131 1.4705
R12466 a_5396_9163.n168 a_5396_9163.t90 1.4705
R12467 a_5396_9163.n168 a_5396_9163.t171 1.4705
R12468 a_5396_9163.n169 a_5396_9163.t127 1.4705
R12469 a_5396_9163.n169 a_5396_9163.t121 1.4705
R12470 a_5396_9163.n172 a_5396_9163.t129 1.4705
R12471 a_5396_9163.n172 a_5396_9163.t130 1.4705
R12472 a_5396_9163.n173 a_5396_9163.t140 1.4705
R12473 a_5396_9163.n173 a_5396_9163.t117 1.4705
R12474 a_5396_9163.n176 a_5396_9163.t88 1.4705
R12475 a_5396_9163.n176 a_5396_9163.t123 1.4705
R12476 a_5396_9163.n177 a_5396_9163.t89 1.4705
R12477 a_5396_9163.n177 a_5396_9163.t108 1.4705
R12478 a_5396_9163.n161 a_5396_9163.t100 1.4705
R12479 a_5396_9163.n161 a_5396_9163.t132 1.4705
R12480 a_5396_9163.n162 a_5396_9163.t101 1.4705
R12481 a_5396_9163.n162 a_5396_9163.t134 1.4705
R12482 a_5396_9163.n157 a_5396_9163.t111 1.4705
R12483 a_5396_9163.n157 a_5396_9163.t156 1.4705
R12484 a_5396_9163.n158 a_5396_9163.t116 1.4705
R12485 a_5396_9163.n158 a_5396_9163.t142 1.4705
R12486 a_5396_9163.n153 a_5396_9163.t144 1.4705
R12487 a_5396_9163.n153 a_5396_9163.t151 1.4705
R12488 a_5396_9163.n154 a_5396_9163.t152 1.4705
R12489 a_5396_9163.n154 a_5396_9163.t96 1.4705
R12490 a_5396_9163.n149 a_5396_9163.t146 1.4705
R12491 a_5396_9163.n149 a_5396_9163.t126 1.4705
R12492 a_5396_9163.n150 a_5396_9163.t147 1.4705
R12493 a_5396_9163.n150 a_5396_9163.t172 1.4705
R12494 a_5396_9163.n100 a_5396_9163.t163 1.4705
R12495 a_5396_9163.n100 a_5396_9163.t159 1.4705
R12496 a_5396_9163.n101 a_5396_9163.t162 1.4705
R12497 a_5396_9163.n101 a_5396_9163.t155 1.4705
R12498 a_5396_9163.n103 a_5396_9163.t107 1.4705
R12499 a_5396_9163.n103 a_5396_9163.t125 1.4705
R12500 a_5396_9163.n104 a_5396_9163.t106 1.4705
R12501 a_5396_9163.n104 a_5396_9163.t124 1.4705
R12502 a_5396_9163.n107 a_5396_9163.t154 1.4705
R12503 a_5396_9163.n107 a_5396_9163.t149 1.4705
R12504 a_5396_9163.n108 a_5396_9163.t153 1.4705
R12505 a_5396_9163.n108 a_5396_9163.t148 1.4705
R12506 a_5396_9163.n111 a_5396_9163.t143 1.4705
R12507 a_5396_9163.n111 a_5396_9163.t93 1.4705
R12508 a_5396_9163.n112 a_5396_9163.t157 1.4705
R12509 a_5396_9163.n112 a_5396_9163.t141 1.4705
R12510 a_5396_9163.n120 a_5396_9163.t114 1.4705
R12511 a_5396_9163.n120 a_5396_9163.t139 1.4705
R12512 a_5396_9163.n121 a_5396_9163.t165 1.4705
R12513 a_5396_9163.n121 a_5396_9163.t138 1.4705
R12514 a_5396_9163.n124 a_5396_9163.t175 1.4705
R12515 a_5396_9163.n124 a_5396_9163.t99 1.4705
R12516 a_5396_9163.n125 a_5396_9163.t174 1.4705
R12517 a_5396_9163.n125 a_5396_9163.t98 1.4705
R12518 a_5396_9163.n128 a_5396_9163.t122 1.4705
R12519 a_5396_9163.n128 a_5396_9163.t135 1.4705
R12520 a_5396_9163.n129 a_5396_9163.t105 1.4705
R12521 a_5396_9163.n129 a_5396_9163.t133 1.4705
R12522 a_5396_9163.n132 a_5396_9163.t91 1.4705
R12523 a_5396_9163.n132 a_5396_9163.t110 1.4705
R12524 a_5396_9163.n133 a_5396_9163.t166 1.4705
R12525 a_5396_9163.n133 a_5396_9163.t160 1.4705
R12526 a_5396_9163.n97 a_5396_9163.t97 1.4705
R12527 a_5396_9163.n97 a_5396_9163.t169 1.4705
R12528 a_5396_9163.n185 a_5396_9163.t103 1.4705
R12529 a_5396_9163.n185 a_5396_9163.t119 1.4705
R12530 a_5396_9163.n146 a_5396_9163.t150 1.4705
R12531 a_5396_9163.n146 a_5396_9163.t167 1.4705
R12532 a_5396_9163.n145 a_5396_9163.t92 1.4705
R12533 a_5396_9163.n145 a_5396_9163.t158 1.4705
R12534 a_5396_9163.n137 a_5396_9163.t137 1.4705
R12535 a_5396_9163.n137 a_5396_9163.t128 1.4705
R12536 a_5396_9163.n141 a_5396_9163.t170 1.4705
R12537 a_5396_9163.n141 a_5396_9163.t164 1.4705
R12538 a_5396_9163.n16 a_5396_9163.n15 1.46537
R12539 a_5396_9163.n18 a_5396_9163.n17 1.46537
R12540 a_5396_9163.n22 a_5396_9163.n21 1.46537
R12541 a_5396_9163.n83 a_5396_9163.n82 1.46537
R12542 a_5396_9163.n85 a_5396_9163.n84 1.46537
R12543 a_5396_9163.n89 a_5396_9163.n88 1.46537
R12544 a_5396_9163.n91 a_5396_9163.n90 1.46537
R12545 a_5396_9163.n81 a_5396_9163.n80 1.46537
R12546 a_5396_9163.n60 a_5396_9163.n59 1.46537
R12547 a_5396_9163.n62 a_5396_9163.n61 1.46537
R12548 a_5396_9163.n55 a_5396_9163.n54 1.46537
R12549 a_5396_9163.n51 a_5396_9163.n50 1.46537
R12550 a_5396_9163.n49 a_5396_9163.n48 1.46537
R12551 a_5396_9163.n47 a_5396_9163.n46 1.46537
R12552 a_5396_9163.n43 a_5396_9163.n42 1.46537
R12553 a_5396_9163.n38 a_5396_9163.n37 1.46537
R12554 a_5396_9163.n171 a_5396_9163.n170 1.46537
R12555 a_5396_9163.n175 a_5396_9163.n174 1.46537
R12556 a_5396_9163.n179 a_5396_9163.n178 1.46537
R12557 a_5396_9163.n164 a_5396_9163.n163 1.46537
R12558 a_5396_9163.n160 a_5396_9163.n159 1.46537
R12559 a_5396_9163.n156 a_5396_9163.n155 1.46537
R12560 a_5396_9163.n152 a_5396_9163.n151 1.46537
R12561 a_5396_9163.n106 a_5396_9163.n105 1.46537
R12562 a_5396_9163.n110 a_5396_9163.n109 1.46537
R12563 a_5396_9163.n114 a_5396_9163.n113 1.46537
R12564 a_5396_9163.n123 a_5396_9163.n122 1.46537
R12565 a_5396_9163.n127 a_5396_9163.n126 1.46537
R12566 a_5396_9163.n131 a_5396_9163.n130 1.46537
R12567 a_5396_9163.n135 a_5396_9163.n134 1.46537
R12568 a_5396_9163.n197 a_5396_9163.n196 1.46535
R12569 a_5396_9163.n93 a_5396_9163.n92 1.46535
R12570 a_5396_9163.n64 a_5396_9163.n63 1.46535
R12571 a_5396_9163.n41 a_5396_9163.n40 1.46535
R12572 a_5396_9163.n30 a_5396_9163.n28 1.27228
R12573 a_5396_9163.n47 a_5396_9163.n43 1.27228
R12574 a_5396_9163.n49 a_5396_9163.n47 1.27228
R12575 a_5396_9163.n55 a_5396_9163.n51 1.27228
R12576 a_5396_9163.n62 a_5396_9163.n60 1.27228
R12577 a_5396_9163.n75 a_5396_9163.n74 1.27228
R12578 a_5396_9163.n91 a_5396_9163.n89 1.27228
R12579 a_5396_9163.n89 a_5396_9163.n85 1.27228
R12580 a_5396_9163.n83 a_5396_9163.n22 1.27228
R12581 a_5396_9163.n18 a_5396_9163.n16 1.27228
R12582 a_5396_9163.n156 a_5396_9163.n152 1.27228
R12583 a_5396_9163.n164 a_5396_9163.n160 1.27228
R12584 a_5396_9163.n179 a_5396_9163.n175 1.27228
R12585 a_5396_9163.n135 a_5396_9163.n131 1.27228
R12586 a_5396_9163.n127 a_5396_9163.n123 1.27228
R12587 a_5396_9163.n114 a_5396_9163.n110 1.27228
R12588 a_5396_9163.n186 a_5396_9163.n184 1.27228
R12589 a_5396_9163.n142 a_5396_9163.n140 1.27228
R12590 a_5396_9163.n182 a_5396_9163.n24 1.25341
R12591 a_5396_9163.n189 a_5396_9163.n188 1.23151
R12592 a_5396_9163.n33 a_5396_9163.n32 1.01873
R12593 a_5396_9163.n72 a_5396_9163.n71 1.01873
R12594 a_5396_9163.n69 a_5396_9163.n25 0.778574
R12595 a_5396_9163.n189 a_5396_9163.n95 0.778574
R12596 a_5396_9163.n67 a_5396_9163.n66 0.778574
R12597 a_5396_9163.n194 a_5396_9163.n193 0.778574
R12598 a_5396_9163.n95 a_5396_9163.n76 0.738439
R12599 a_5396_9163.n194 a_5396_9163.n23 0.738439
R12600 a_5396_9163.n187 a_5396_9163.n96 0.737223
R12601 a_5396_9163.n143 a_5396_9163.n136 0.737223
R12602 a_5396_9163.n182 a_5396_9163.n181 0.737223
R12603 a_5396_9163.n118 a_5396_9163.n99 0.737223
R12604 a_5396_9163.n144 a_5396_9163.n143 0.725061
R12605 a_5396_9163.n148 a_5396_9163.n99 0.725061
R12606 a_5396_9163.n41 a_5396_9163.n39 0.699581
R12607 a_5396_9163.n65 a_5396_9163.n64 0.699581
R12608 a_5396_9163.n94 a_5396_9163.n93 0.699581
R12609 a_5396_9163.n196 a_5396_9163.n195 0.699581
R12610 a_5396_9163.n144 a_5396_9163.n96 0.585196
R12611 a_5396_9163.n181 a_5396_9163.n148 0.585196
R12612 a_5396_9163.n39 a_5396_9163.n38 0.557791
R12613 a_5396_9163.n65 a_5396_9163.n55 0.557791
R12614 a_5396_9163.n94 a_5396_9163.n81 0.557791
R12615 a_5396_9163.n195 a_5396_9163.n22 0.557791
R12616 a_5396_9163.n76 a_5396_9163.n69 0.530466
R12617 a_5396_9163.n67 a_5396_9163.n23 0.530466
R12618 a_5396_9163.n180 a_5396_9163.n179 0.150184
R12619 a_5396_9163.n119 a_5396_9163.n114 0.150184
R12620 a_5396_9163.n1 a_5396_9163.n2 1.27228
R12621 a_5396_9163.n68 a_5396_9163.n1 7.30549
R12622 a_5396_9163.t71 a_5396_9163.n0 6.96214
R12623 a_5396_9163.n4 a_5396_9163.n5 1.27228
R12624 a_5396_9163.n192 a_5396_9163.n4 7.30549
R12625 a_5396_9163.t58 a_5396_9163.n3 6.96214
R12626 a_5396_9163.n10 a_5396_9163.n11 1.26457
R12627 a_5396_9163.n147 a_5396_9163.n10 6.59229
R12628 a_5396_9163.n146 a_5396_9163.n9 5.10549
R12629 a_5396_9163.n7 a_5396_9163.n8 1.26457
R12630 a_5396_9163.n117 a_5396_9163.n7 6.59229
R12631 a_5396_9163.n116 a_5396_9163.n6 5.10549
R12632 VOUT.n24 VOUT.n17 7.94229
R12633 VOUT.n77 VOUT.n75 7.94229
R12634 VOUT.n72 VOUT.n65 7.169
R12635 VOUT.n138 VOUT.n137 7.169
R12636 VOUT.n117 VOUT.t104 6.96668
R12637 VOUT.n8 VOUT.t49 6.82564
R12638 VOUT.n69 VOUT.t71 6.82564
R12639 VOUT.n133 VOUT.t93 5.85326
R12640 VOUT.n133 VOUT.n132 5.84661
R12641 VOUT.n16 VOUT.t23 5.69423
R12642 VOUT.n25 VOUT.t65 5.69423
R12643 VOUT.n14 VOUT.t87 5.69423
R12644 VOUT.n78 VOUT.t10 5.69423
R12645 VOUT.n16 VOUT.n15 5.49558
R12646 VOUT.n14 VOUT.n13 5.49558
R12647 VOUT.n10 VOUT.n9 4.61332
R12648 VOUT.n140 VOUT.n139 4.61332
R12649 VOUT.n71 VOUT.n70 4.61332
R12650 VOUT.n64 VOUT.n62 4.61332
R12651 VOUT.n60 VOUT.n57 4.61332
R12652 VOUT.n119 VOUT.n118 4.61332
R12653 VOUT.n2 VOUT.n1 4.61332
R12654 VOUT.n9 VOUT.n8 4.60571
R12655 VOUT.n139 VOUT.n138 4.60571
R12656 VOUT.n70 VOUT.n69 4.60571
R12657 VOUT.n65 VOUT.n64 4.60571
R12658 VOUT.n61 VOUT.n60 4.60571
R12659 VOUT.n118 VOUT.n117 4.60571
R12660 VOUT.n141 VOUT.n1 4.60571
R12661 VOUT.n59 VOUT.n56 4.5005
R12662 VOUT.n63 VOUT.n55 4.5005
R12663 VOUT.n68 VOUT.n66 4.5005
R12664 VOUT.n116 VOUT.n114 4.5005
R12665 VOUT.n4 VOUT.n3 4.5005
R12666 VOUT.n7 VOUT.n5 4.5005
R12667 VOUT.n143 VOUT.n142 4.5005
R12668 VOUT.n4 VOUT.t64 4.22462
R12669 VOUT.n63 VOUT.t30 4.22462
R12670 VOUT.n24 VOUT.n23 4.22423
R12671 VOUT.n77 VOUT.n76 4.22423
R12672 VOUT.n126 VOUT.t91 4.21195
R12673 VOUT.n128 VOUT.t94 4.21195
R12674 VOUT.n44 VOUT.t55 4.05054
R12675 VOUT.n49 VOUT.t75 4.05054
R12676 VOUT.n51 VOUT.t57 4.05054
R12677 VOUT.n38 VOUT.t41 4.05054
R12678 VOUT.n36 VOUT.t16 4.05054
R12679 VOUT.n30 VOUT.t56 4.05054
R12680 VOUT.n28 VOUT.t22 4.05054
R12681 VOUT.n18 VOUT.t81 4.05054
R12682 VOUT.n85 VOUT.t29 4.05054
R12683 VOUT.n90 VOUT.t46 4.05054
R12684 VOUT.n92 VOUT.t4 4.05054
R12685 VOUT.n99 VOUT.t83 4.05054
R12686 VOUT.n101 VOUT.t42 4.05054
R12687 VOUT.n107 VOUT.t38 4.05054
R12688 VOUT.n109 VOUT.t15 4.05054
R12689 VOUT.n80 VOUT.t70 4.05054
R12690 VOUT.n126 VOUT.t98 4.03668
R12691 VOUT.n128 VOUT.t101 4.03668
R12692 VOUT.n44 VOUT.t51 3.87765
R12693 VOUT.n49 VOUT.t72 3.87765
R12694 VOUT.n51 VOUT.t54 3.87765
R12695 VOUT.n38 VOUT.t40 3.87765
R12696 VOUT.n36 VOUT.t14 3.87765
R12697 VOUT.n30 VOUT.t53 3.87765
R12698 VOUT.n28 VOUT.t21 3.87765
R12699 VOUT.n18 VOUT.t80 3.87765
R12700 VOUT.n85 VOUT.t31 3.87765
R12701 VOUT.n90 VOUT.t47 3.87765
R12702 VOUT.n92 VOUT.t5 3.87765
R12703 VOUT.n99 VOUT.t85 3.87765
R12704 VOUT.n101 VOUT.t43 3.87765
R12705 VOUT.n107 VOUT.t39 3.87765
R12706 VOUT.n109 VOUT.t17 3.87765
R12707 VOUT.n80 VOUT.t73 3.87765
R12708 VOUT.n131 VOUT.n119 3.81532
R12709 VOUT.n136 VOUT.n135 3.544
R12710 VOUT.n135 VOUT.n113 3.48165
R12711 VOUT.n26 VOUT.n25 3.25667
R12712 VOUT.n116 VOUT.n115 3.12366
R12713 VOUT.n57 VOUT.n12 3.01925
R12714 VOUT.n113 VOUT.n2 3.01925
R12715 VOUT.n125 VOUT.n124 2.95195
R12716 VOUT.n122 VOUT.n121 2.95195
R12717 VOUT.n125 VOUT.n123 2.77668
R12718 VOUT.n122 VOUT.n120 2.77668
R12719 VOUT.n7 VOUT.n6 2.75462
R12720 VOUT.n68 VOUT.n67 2.75462
R12721 VOUT.n59 VOUT.n58 2.75462
R12722 VOUT.n22 VOUT.n18 2.73714
R12723 VOUT.n84 VOUT.n80 2.73714
R12724 VOUT.n48 VOUT.n44 2.73672
R12725 VOUT.n89 VOUT.n85 2.73672
R12726 VOUT.n127 VOUT.n125 2.71872
R12727 VOUT.n39 VOUT.n37 2.60203
R12728 VOUT.n102 VOUT.n100 2.60203
R12729 VOUT.n47 VOUT.n46 2.58054
R12730 VOUT.n42 VOUT.n41 2.58054
R12731 VOUT.n34 VOUT.n33 2.58054
R12732 VOUT.n21 VOUT.n20 2.58054
R12733 VOUT.n88 VOUT.n87 2.58054
R12734 VOUT.n97 VOUT.n96 2.58054
R12735 VOUT.n105 VOUT.n104 2.58054
R12736 VOUT.n83 VOUT.n82 2.58054
R12737 VOUT.n129 VOUT.n127 2.56118
R12738 VOUT.n134 VOUT.n133 2.54573
R12739 VOUT.n31 VOUT.n29 2.53418
R12740 VOUT.n52 VOUT.n50 2.53418
R12741 VOUT.n110 VOUT.n108 2.53418
R12742 VOUT.n93 VOUT.n91 2.53418
R12743 VOUT.n79 VOUT.n78 2.51873
R12744 VOUT.n47 VOUT.n45 2.40765
R12745 VOUT.n42 VOUT.n40 2.40765
R12746 VOUT.n34 VOUT.n32 2.40765
R12747 VOUT.n21 VOUT.n19 2.40765
R12748 VOUT.n88 VOUT.n86 2.40765
R12749 VOUT.n97 VOUT.n95 2.40765
R12750 VOUT.n105 VOUT.n103 2.40765
R12751 VOUT.n83 VOUT.n81 2.40765
R12752 VOUT.n54 VOUT.n17 2.23844
R12753 VOUT VOUT.n0 2.05949
R12754 VOUT.n130 VOUT.n122 2.00466
R12755 VOUT.n72 VOUT.n71 1.51925
R12756 VOUT.n137 VOUT.n10 1.51925
R12757 VOUT.n112 VOUT.n111 1.5005
R12758 VOUT.n27 VOUT.n26 1.5005
R12759 VOUT.n131 VOUT.n130 1.5005
R12760 VOUT.n94 VOUT.n11 1.5005
R12761 VOUT.n75 VOUT.n74 1.5005
R12762 VOUT.n73 VOUT.n72 1.5005
R12763 VOUT.n54 VOUT.n53 1.5005
R12764 VOUT.n137 VOUT.n136 1.5005
R12765 VOUT.n0 VOUT.t25 1.4705
R12766 VOUT.n0 VOUT.t86 1.4705
R12767 VOUT.n6 VOUT.t12 1.4705
R12768 VOUT.n6 VOUT.t69 1.4705
R12769 VOUT.n15 VOUT.t45 1.4705
R12770 VOUT.n15 VOUT.t44 1.4705
R12771 VOUT.n23 VOUT.t3 1.4705
R12772 VOUT.n23 VOUT.t2 1.4705
R12773 VOUT.n45 VOUT.t11 1.4705
R12774 VOUT.n45 VOUT.t6 1.4705
R12775 VOUT.n46 VOUT.t13 1.4705
R12776 VOUT.n46 VOUT.t7 1.4705
R12777 VOUT.n40 VOUT.t35 1.4705
R12778 VOUT.n40 VOUT.t59 1.4705
R12779 VOUT.n41 VOUT.t36 1.4705
R12780 VOUT.n41 VOUT.t60 1.4705
R12781 VOUT.n32 VOUT.t82 1.4705
R12782 VOUT.n32 VOUT.t78 1.4705
R12783 VOUT.n33 VOUT.t84 1.4705
R12784 VOUT.n33 VOUT.t79 1.4705
R12785 VOUT.n19 VOUT.t74 1.4705
R12786 VOUT.n19 VOUT.t24 1.4705
R12787 VOUT.n20 VOUT.t76 1.4705
R12788 VOUT.n20 VOUT.t26 1.4705
R12789 VOUT.n67 VOUT.t77 1.4705
R12790 VOUT.n67 VOUT.t20 1.4705
R12791 VOUT.n58 VOUT.t32 1.4705
R12792 VOUT.n58 VOUT.t62 1.4705
R12793 VOUT.n13 VOUT.t58 1.4705
R12794 VOUT.n13 VOUT.t37 1.4705
R12795 VOUT.n76 VOUT.t66 1.4705
R12796 VOUT.n76 VOUT.t48 1.4705
R12797 VOUT.n86 VOUT.t19 1.4705
R12798 VOUT.n86 VOUT.t1 1.4705
R12799 VOUT.n87 VOUT.t18 1.4705
R12800 VOUT.n87 VOUT.t0 1.4705
R12801 VOUT.n95 VOUT.t63 1.4705
R12802 VOUT.n95 VOUT.t28 1.4705
R12803 VOUT.n96 VOUT.t61 1.4705
R12804 VOUT.n96 VOUT.t27 1.4705
R12805 VOUT.n103 VOUT.t9 1.4705
R12806 VOUT.n103 VOUT.t68 1.4705
R12807 VOUT.n104 VOUT.t8 1.4705
R12808 VOUT.n104 VOUT.t67 1.4705
R12809 VOUT.n81 VOUT.t52 1.4705
R12810 VOUT.n81 VOUT.t34 1.4705
R12811 VOUT.n82 VOUT.t50 1.4705
R12812 VOUT.n82 VOUT.t33 1.4705
R12813 VOUT.n48 VOUT.n47 1.46537
R12814 VOUT.n50 VOUT.n49 1.46537
R12815 VOUT.n43 VOUT.n42 1.46537
R12816 VOUT.n39 VOUT.n38 1.46537
R12817 VOUT.n37 VOUT.n36 1.46537
R12818 VOUT.n35 VOUT.n34 1.46537
R12819 VOUT.n31 VOUT.n30 1.46537
R12820 VOUT.n22 VOUT.n21 1.46537
R12821 VOUT.n89 VOUT.n88 1.46537
R12822 VOUT.n91 VOUT.n90 1.46537
R12823 VOUT.n98 VOUT.n97 1.46537
R12824 VOUT.n100 VOUT.n99 1.46537
R12825 VOUT.n102 VOUT.n101 1.46537
R12826 VOUT.n106 VOUT.n105 1.46537
R12827 VOUT.n108 VOUT.n107 1.46537
R12828 VOUT.n84 VOUT.n83 1.46537
R12829 VOUT.n127 VOUT.n126 1.46537
R12830 VOUT.n52 VOUT.n51 1.46535
R12831 VOUT.n29 VOUT.n28 1.46535
R12832 VOUT.n93 VOUT.n92 1.46535
R12833 VOUT.n110 VOUT.n109 1.46535
R12834 VOUT.n129 VOUT.n128 1.46535
R12835 VOUT.n25 VOUT.n24 1.27228
R12836 VOUT.n35 VOUT.n31 1.27228
R12837 VOUT.n37 VOUT.n35 1.27228
R12838 VOUT.n43 VOUT.n39 1.27228
R12839 VOUT.n50 VOUT.n48 1.27228
R12840 VOUT.n78 VOUT.n77 1.27228
R12841 VOUT.n108 VOUT.n106 1.27228
R12842 VOUT.n106 VOUT.n102 1.27228
R12843 VOUT.n100 VOUT.n98 1.27228
R12844 VOUT.n91 VOUT.n89 1.27228
R12845 VOUT.n132 VOUT.t99 1.2605
R12846 VOUT.n132 VOUT.t92 1.2605
R12847 VOUT.n123 VOUT.t103 1.2605
R12848 VOUT.n123 VOUT.t97 1.2605
R12849 VOUT.n124 VOUT.t96 1.2605
R12850 VOUT.n124 VOUT.t90 1.2605
R12851 VOUT.n120 VOUT.t102 1.2605
R12852 VOUT.n120 VOUT.t88 1.2605
R12853 VOUT.n121 VOUT.t95 1.2605
R12854 VOUT.n121 VOUT.t100 1.2605
R12855 VOUT.n115 VOUT.t105 1.2605
R12856 VOUT.n115 VOUT.t89 1.2605
R12857 VOUT.n135 VOUT.n134 1.25797
R12858 VOUT.n17 VOUT.n16 1.01873
R12859 VOUT.n75 VOUT.n14 1.01873
R12860 VOUT.n62 VOUT.n61 0.9995
R12861 VOUT.n141 VOUT.n140 0.9995
R12862 VOUT.n26 VOUT.n12 0.778574
R12863 VOUT.n113 VOUT.n112 0.778574
R12864 VOUT.n73 VOUT.n54 0.778574
R12865 VOUT.n136 VOUT.n11 0.778574
R12866 VOUT.n112 VOUT.n79 0.738439
R12867 VOUT.n134 VOUT.n131 0.738439
R12868 VOUT.n74 VOUT.n11 0.738439
R12869 VOUT.n29 VOUT.n27 0.699581
R12870 VOUT.n53 VOUT.n52 0.699581
R12871 VOUT.n111 VOUT.n110 0.699581
R12872 VOUT.n94 VOUT.n93 0.699581
R12873 VOUT.n130 VOUT.n129 0.699581
R12874 VOUT VOUT.n143 0.695632
R12875 VOUT.n27 VOUT.n22 0.557791
R12876 VOUT.n53 VOUT.n43 0.557791
R12877 VOUT.n111 VOUT.n84 0.557791
R12878 VOUT.n98 VOUT.n94 0.557791
R12879 VOUT.n79 VOUT.n12 0.530466
R12880 VOUT.n74 VOUT.n73 0.530466
R12881 VOUT.n57 VOUT.n56 0.14
R12882 VOUT.n61 VOUT.n56 0.14
R12883 VOUT.n62 VOUT.n55 0.14
R12884 VOUT.n65 VOUT.n55 0.14
R12885 VOUT.n71 VOUT.n66 0.14
R12886 VOUT.n69 VOUT.n66 0.14
R12887 VOUT.n119 VOUT.n114 0.14
R12888 VOUT.n117 VOUT.n114 0.14
R12889 VOUT.n142 VOUT.n2 0.14
R12890 VOUT.n142 VOUT.n141 0.14
R12891 VOUT.n140 VOUT.n3 0.14
R12892 VOUT.n138 VOUT.n3 0.14
R12893 VOUT.n10 VOUT.n5 0.14
R12894 VOUT.n8 VOUT.n5 0.14
R12895 VOUT.n9 VOUT.n7 0.00168421
R12896 VOUT.n139 VOUT.n4 0.00168421
R12897 VOUT.n70 VOUT.n68 0.00168421
R12898 VOUT.n64 VOUT.n63 0.00168421
R12899 VOUT.n60 VOUT.n59 0.00168421
R12900 VOUT.n118 VOUT.n116 0.00168421
R12901 VOUT.n143 VOUT.n1 0.00168421
R12902 a_n11737_n14973.n334 a_n11737_n14973.t4 10.621
R12903 a_n11737_n14973.n330 a_n11737_n14973.t35 10.621
R12904 a_n11737_n14973.n340 a_n11737_n14973.n328 10.3121
R12905 a_n11737_n14973.n336 a_n11737_n14973.t77 10.3044
R12906 a_n11737_n14973.n332 a_n11737_n14973.t6 10.3044
R12907 a_n11737_n14973.n335 a_n11737_n14973.t95 9.9994
R12908 a_n11737_n14973.n331 a_n11737_n14973.t2 9.9994
R12909 a_n11737_n14973.n334 a_n11737_n14973.t0 9.999
R12910 a_n11737_n14973.n330 a_n11737_n14973.t48 9.999
R12911 a_n11737_n14973.n226 a_n11737_n14973.t54 8.33806
R12912 a_n11737_n14973.n321 a_n11737_n14973.t93 8.3366
R12913 a_n11737_n14973.n280 a_n11737_n14973.t76 8.26493
R12914 a_n11737_n14973.n96 a_n11737_n14973.t69 8.35715
R12915 a_n11737_n14973.n43 a_n11737_n14973.t99 8.06917
R12916 a_n11737_n14973.n55 a_n11737_n14973.t67 8.06917
R12917 a_n11737_n14973.n122 a_n11737_n14973.t90 8.06917
R12918 a_n11737_n14973.n31 a_n11737_n14973.t75 8.06917
R12919 a_n11737_n14973.n132 a_n11737_n14973.t104 8.06917
R12920 a_n11737_n14973.n50 a_n11737_n14973.t55 8.06917
R12921 a_n11737_n14973.n57 a_n11737_n14973.t31 8.06917
R12922 a_n11737_n14973.n17 a_n11737_n14973.t44 8.06917
R12923 a_n11737_n14973.n78 a_n11737_n14973.t33 8.06917
R12924 a_n11737_n14973.n28 a_n11737_n14973.t84 8.06917
R12925 a_n11737_n14973.n133 a_n11737_n14973.t32 8.06917
R12926 a_n11737_n14973.n9 a_n11737_n14973.t47 8.06917
R12927 a_n11737_n14973.n8 a_n11737_n14973.t34 8.06917
R12928 a_n11737_n14973.n172 a_n11737_n14973.t45 8.06917
R12929 a_n11737_n14973.n6 a_n11737_n14973.t79 8.06917
R12930 a_n11737_n14973.n5 a_n11737_n14973.t57 8.06917
R12931 a_n11737_n14973.n177 a_n11737_n14973.t78 8.06917
R12932 a_n11737_n14973.n40 a_n11737_n14973.t66 8.06917
R12933 a_n11737_n14973.n93 a_n11737_n14973.t74 8.06917
R12934 a_n11737_n14973.n75 a_n11737_n14973.t49 8.06917
R12935 a_n11737_n14973.n61 a_n11737_n14973.t73 8.06917
R12936 a_n11737_n14973.n34 a_n11737_n14973.t30 8.06917
R12937 a_n11737_n14973.n90 a_n11737_n14973.t80 8.06917
R12938 a_n11737_n14973.n2 a_n11737_n14973.t100 8.06917
R12939 a_n11737_n14973.n86 a_n11737_n14973.t82 8.06917
R12940 a_n11737_n14973.n71 a_n11737_n14973.t53 8.06917
R12941 a_n11737_n14973.n65 a_n11737_n14973.t81 8.06917
R12942 a_n11737_n14973.n125 a_n11737_n14973.t64 8.06917
R12943 a_n11737_n14973.n23 a_n11737_n14973.t50 8.06917
R12944 a_n11737_n14973.n165 a_n11737_n14973.t63 8.06917
R12945 a_n11737_n14973.n128 a_n11737_n14973.t102 8.06917
R12946 a_n11737_n14973.n20 a_n11737_n14973.t86 8.06917
R12947 a_n11737_n14973.n154 a_n11737_n14973.t101 8.06917
R12948 a_n11737_n14973.n82 a_n11737_n14973.t41 8.06917
R12949 a_n11737_n14973.n68 a_n11737_n14973.t58 8.06917
R12950 a_n11737_n14973.n108 a_n11737_n14973.t103 8.06917
R12951 a_n11737_n14973.n97 a_n11737_n14973.t70 8.06917
R12952 a_n11737_n14973.n261 a_n11737_n14973.t91 8.06917
R12953 a_n11737_n14973.n250 a_n11737_n14973.t83 8.06917
R12954 a_n11737_n14973.n249 a_n11737_n14973.t59 8.06917
R12955 a_n11737_n14973.n248 a_n11737_n14973.t85 8.06917
R12956 a_n11737_n14973.n95 a_n11737_n14973.t42 8.06917
R12957 a_n11737_n14973.n241 a_n11737_n14973.t68 8.06917
R12958 a_n11737_n14973.n112 a_n11737_n14973.t60 8.06917
R12959 a_n11737_n14973.n227 a_n11737_n14973.t40 8.06917
R12960 a_n11737_n14973.n233 a_n11737_n14973.t36 8.06917
R12961 a_n11737_n14973.n234 a_n11737_n14973.t94 8.06917
R12962 a_n11737_n14973.n235 a_n11737_n14973.t37 8.06917
R12963 a_n11737_n14973.n109 a_n11737_n14973.t72 8.06917
R12964 a_n11737_n14973.n100 a_n11737_n14973.t46 8.06917
R12965 a_n11737_n14973.n269 a_n11737_n14973.t71 8.06917
R12966 a_n11737_n14973.n320 a_n11737_n14973.t61 8.06917
R12967 a_n11737_n14973.n118 a_n11737_n14973.t92 8.06917
R12968 a_n11737_n14973.n318 a_n11737_n14973.t52 8.06917
R12969 a_n11737_n14973.n317 a_n11737_n14973.t38 8.06917
R12970 a_n11737_n14973.n316 a_n11737_n14973.t51 8.06917
R12971 a_n11737_n14973.n314 a_n11737_n14973.t43 8.06917
R12972 a_n11737_n14973.n307 a_n11737_n14973.t96 8.06917
R12973 a_n11737_n14973.n115 a_n11737_n14973.t39 8.06917
R12974 a_n11737_n14973.n302 a_n11737_n14973.t98 8.06917
R12975 a_n11737_n14973.n101 a_n11737_n14973.t65 8.06917
R12976 a_n11737_n14973.n119 a_n11737_n14973.t97 8.06917
R12977 a_n11737_n14973.n291 a_n11737_n14973.t88 8.06917
R12978 a_n11737_n14973.n290 a_n11737_n14973.t62 8.06917
R12979 a_n11737_n14973.n289 a_n11737_n14973.t87 8.06917
R12980 a_n11737_n14973.n276 a_n11737_n14973.t89 8.06917
R12981 a_n11737_n14973.n279 a_n11737_n14973.t56 8.06917
R12982 a_n11737_n14973.t29 a_n11737_n14973.n359 6.49245
R12983 a_n11737_n14973.n143 a_n11737_n14973.t15 6.49245
R12984 a_n11737_n14973.n140 a_n11737_n14973.t23 6.50349
R12985 a_n11737_n14973.n338 a_n11737_n14973.t5 5.70664
R12986 a_n11737_n14973.n329 a_n11737_n14973.t7 5.23357
R12987 a_n11737_n14973.n144 a_n11737_n14973.t18 5.22068
R12988 a_n11737_n14973.n329 a_n11737_n14973.t3 5.15078
R12989 a_n11737_n14973.n338 a_n11737_n14973.t1 4.6582
R12990 a_n11737_n14973.n84 a_n11737_n14973.n69 2.0194
R12991 a_n11737_n14973.n180 a_n11737_n14973.n123 2.42484
R12992 a_n11737_n14973.n123 a_n11737_n14973.n179 2.4256
R12993 a_n11737_n14973.n110 a_n11737_n14973.n109 2.25048
R12994 a_n11737_n14973.n115 a_n11737_n14973.n113 2.25048
R12995 a_n11737_n14973.n136 a_n11737_n14973.n342 3.76239
R12996 a_n11737_n14973.n137 a_n11737_n14973.t14 5.23239
R12997 a_n11737_n14973.n349 a_n11737_n14973.n348 4.60825
R12998 a_n11737_n14973.n345 a_n11737_n14973.n140 3.76239
R12999 a_n11737_n14973.n10 a_n11737_n14973.n9 1.44552
R13000 a_n11737_n14973.n7 a_n11737_n14973.n6 1.44552
R13001 a_n11737_n14973.n126 a_n11737_n14973.n125 2.22591
R13002 a_n11737_n14973.n129 a_n11737_n14973.n128 2.22591
R13003 a_n11737_n14973.n85 a_n11737_n14973.n161 4.51491
R13004 a_n11737_n14973.n218 a_n11737_n14973.n217 4.51075
R13005 a_n11737_n14973.n62 a_n11737_n14973.n61 2.21906
R13006 a_n11737_n14973.n66 a_n11737_n14973.n65 2.21906
R13007 a_n11737_n14973.n34 a_n11737_n14973.n35 2.21826
R13008 a_n11737_n14973.n40 a_n11737_n14973.n39 2.21826
R13009 a_n11737_n14973.n348 a_n11737_n14973.n341 4.50168
R13010 a_n11737_n14973.n347 a_n11737_n14973.n346 4.5005
R13011 a_n11737_n14973.n139 a_n11737_n14973.n138 2.24327
R13012 a_n11737_n14973.n12 a_n11737_n14973.n5 2.21666
R13013 a_n11737_n14973.n11 a_n11737_n14973.n176 4.5005
R13014 a_n11737_n14973.n186 a_n11737_n14973.n185 4.5005
R13015 a_n11737_n14973.n14 a_n11737_n14973.n8 2.21666
R13016 a_n11737_n14973.n13 a_n11737_n14973.n171 4.5005
R13017 a_n11737_n14973.n204 a_n11737_n14973.n203 4.5005
R13018 a_n11737_n14973.n196 a_n11737_n14973.n195 4.5005
R13019 a_n11737_n14973.n78 a_n11737_n14973.n79 2.21666
R13020 a_n11737_n14973.n193 a_n11737_n14973.n27 4.5005
R13021 a_n11737_n14973.n28 a_n11737_n14973.n25 2.21666
R13022 a_n11737_n14973.n26 a_n11737_n14973.n192 4.5005
R13023 a_n11737_n14973.n191 a_n11737_n14973.n133 4.5005
R13024 a_n11737_n14973.n190 a_n11737_n14973.n189 4.5005
R13025 a_n11737_n14973.n51 a_n11737_n14973.n50 2.21666
R13026 a_n11737_n14973.n198 a_n11737_n14973.n49 4.5005
R13027 a_n11737_n14973.n200 a_n11737_n14973.n199 4.5005
R13028 a_n11737_n14973.n58 a_n11737_n14973.n57 2.21666
R13029 a_n11737_n14973.n16 a_n11737_n14973.n173 4.5005
R13030 a_n11737_n14973.n18 a_n11737_n14973.n17 2.21666
R13031 a_n11737_n14973.n0 a_n11737_n14973.n1 0.0657695
R13032 a_n11737_n14973.n30 a_n11737_n14973.n208 4.5005
R13033 a_n11737_n14973.n32 a_n11737_n14973.n31 2.21666
R13034 a_n11737_n14973.n131 a_n11737_n14973.n207 4.5005
R13035 a_n11737_n14973.n132 a_n11737_n14973.n206 4.5005
R13036 a_n11737_n14973.n210 a_n11737_n14973.n205 4.5005
R13037 a_n11737_n14973.n44 a_n11737_n14973.n43 2.21666
R13038 a_n11737_n14973.n42 a_n11737_n14973.n183 4.5005
R13039 a_n11737_n14973.n182 a_n11737_n14973.n54 4.5005
R13040 a_n11737_n14973.n55 a_n11737_n14973.n52 2.21666
R13041 a_n11737_n14973.n53 a_n11737_n14973.n180 4.5005
R13042 a_n11737_n14973.n123 a_n11737_n14973.n122 0.0107891
R13043 a_n11737_n14973.n127 a_n11737_n14973.n160 4.5005
R13044 a_n11737_n14973.n21 a_n11737_n14973.n20 2.21666
R13045 a_n11737_n14973.n19 a_n11737_n14973.n153 4.5005
R13046 a_n11737_n14973.n159 a_n11737_n14973.n158 4.5005
R13047 a_n11737_n14973.n124 a_n11737_n14973.n168 4.5005
R13048 a_n11737_n14973.n24 a_n11737_n14973.n23 2.21666
R13049 a_n11737_n14973.n22 a_n11737_n14973.n164 4.5005
R13050 a_n11737_n14973.n167 a_n11737_n14973.n166 4.5005
R13051 a_n11737_n14973.n65 a_n11737_n14973.n67 2.21666
R13052 a_n11737_n14973.n64 a_n11737_n14973.n107 4.5005
R13053 a_n11737_n14973.n71 a_n11737_n14973.n73 2.21666
R13054 a_n11737_n14973.n70 a_n11737_n14973.n105 4.5005
R13055 a_n11737_n14973.n86 a_n11737_n14973.n88 2.21666
R13056 a_n11737_n14973.n217 a_n11737_n14973.n216 4.5005
R13057 a_n11737_n14973.n2 a_n11737_n14973.n3 2.21666
R13058 a_n11737_n14973.n90 a_n11737_n14973.n92 2.21666
R13059 a_n11737_n14973.n89 a_n11737_n14973.n102 4.5005
R13060 a_n11737_n14973.n162 a_n11737_n14973.n120 4.5005
R13061 a_n11737_n14973.n36 a_n11737_n14973.n34 2.21666
R13062 a_n11737_n14973.n61 a_n11737_n14973.n63 2.21666
R13063 a_n11737_n14973.n60 a_n11737_n14973.n106 4.5005
R13064 a_n11737_n14973.n75 a_n11737_n14973.n77 2.21666
R13065 a_n11737_n14973.n74 a_n11737_n14973.n104 4.5005
R13066 a_n11737_n14973.n68 a_n11737_n14973.n69 0.0231698
R13067 a_n11737_n14973.n82 a_n11737_n14973.n84 2.21666
R13068 a_n11737_n14973.n155 a_n11737_n14973.n81 4.5005
R13069 a_n11737_n14973.n121 a_n11737_n14973.n156 4.5005
R13070 a_n11737_n14973.n41 a_n11737_n14973.n40 2.21666
R13071 a_n11737_n14973.n83 a_n11737_n14973.n82 2.21666
R13072 a_n11737_n14973.n81 a_n11737_n14973.n103 4.5005
R13073 a_n11737_n14973.n38 a_n11737_n14973.n121 4.5005
R13074 a_n11737_n14973.n64 a_n11737_n14973.n221 4.5005
R13075 a_n11737_n14973.n72 a_n11737_n14973.n71 2.21666
R13076 a_n11737_n14973.n70 a_n11737_n14973.n220 4.5005
R13077 a_n11737_n14973.n87 a_n11737_n14973.n86 2.21666
R13078 a_n11737_n14973.n85 a_n11737_n14973.n219 4.5005
R13079 a_n11737_n14973.n2 a_n11737_n14973.n4 2.21666
R13080 a_n11737_n14973.n91 a_n11737_n14973.n90 2.21666
R13081 a_n11737_n14973.n89 a_n11737_n14973.n215 4.5005
R13082 a_n11737_n14973.n214 a_n11737_n14973.n120 4.5005
R13083 a_n11737_n14973.n60 a_n11737_n14973.n170 4.5005
R13084 a_n11737_n14973.n76 a_n11737_n14973.n75 2.21666
R13085 a_n11737_n14973.n74 a_n11737_n14973.n169 4.5005
R13086 a_n11737_n14973.n94 a_n11737_n14973.n93 0.023589
R13087 a_n11737_n14973.n56 a_n11737_n14973.n55 2.21666
R13088 a_n11737_n14973.n181 a_n11737_n14973.n54 4.5005
R13089 a_n11737_n14973.n42 a_n11737_n14973.n178 4.5005
R13090 a_n11737_n14973.n43 a_n11737_n14973.n45 2.21666
R13091 a_n11737_n14973.n53 a_n11737_n14973.n179 4.5005
R13092 a_n11737_n14973.n80 a_n11737_n14973.n78 2.21666
R13093 a_n11737_n14973.n195 a_n11737_n14973.n194 4.5005
R13094 a_n11737_n14973.n189 a_n11737_n14973.n188 4.5005
R13095 a_n11737_n14973.n187 a_n11737_n14973.n133 4.5005
R13096 a_n11737_n14973.n26 a_n11737_n14973.n175 4.5005
R13097 a_n11737_n14973.n29 a_n11737_n14973.n28 2.21666
R13098 a_n11737_n14973.n27 a_n11737_n14973.n174 4.5005
R13099 a_n11737_n14973.n57 a_n11737_n14973.n59 2.21666
R13100 a_n11737_n14973.n201 a_n11737_n14973.n200 4.5005
R13101 a_n11737_n14973.n47 a_n11737_n14973.n49 4.5005
R13102 a_n11737_n14973.n50 a_n11737_n14973.n48 2.21666
R13103 a_n11737_n14973.n17 a_n11737_n14973.n15 2.21666
R13104 a_n11737_n14973.n197 a_n11737_n14973.n16 4.5005
R13105 a_n11737_n14973.n211 a_n11737_n14973.n210 4.5005
R13106 a_n11737_n14973.n132 a_n11737_n14973.n130 4.5005
R13107 a_n11737_n14973.n131 a_n11737_n14973.n209 4.5005
R13108 a_n11737_n14973.n33 a_n11737_n14973.n31 2.21666
R13109 a_n11737_n14973.n30 a_n11737_n14973.n0 0.0743189
R13110 a_n11737_n14973.n301 a_n11737_n14973.n150 4.5005
R13111 a_n11737_n14973.n281 a_n11737_n14973.n278 4.5005
R13112 a_n11737_n14973.n283 a_n11737_n14973.n282 4.5005
R13113 a_n11737_n14973.n284 a_n11737_n14973.n277 4.5005
R13114 a_n11737_n14973.n286 a_n11737_n14973.n285 4.5005
R13115 a_n11737_n14973.n288 a_n11737_n14973.n287 4.5005
R13116 a_n11737_n14973.n293 a_n11737_n14973.n292 4.5005
R13117 a_n11737_n14973.n119 a_n11737_n14973.n294 4.5005
R13118 a_n11737_n14973.n295 a_n11737_n14973.n151 4.5005
R13119 a_n11737_n14973.n297 a_n11737_n14973.n296 4.5005
R13120 a_n11737_n14973.n298 a_n11737_n14973.n101 4.5005
R13121 a_n11737_n14973.n300 a_n11737_n14973.n299 4.5005
R13122 a_n11737_n14973.n304 a_n11737_n14973.n114 4.5005
R13123 a_n11737_n14973.n306 a_n11737_n14973.n305 4.5005
R13124 a_n11737_n14973.n308 a_n11737_n14973.n149 4.5005
R13125 a_n11737_n14973.n310 a_n11737_n14973.n309 4.5005
R13126 a_n11737_n14973.n311 a_n11737_n14973.n148 4.5005
R13127 a_n11737_n14973.n313 a_n11737_n14973.n312 4.5005
R13128 a_n11737_n14973.n315 a_n11737_n14973.n147 4.5005
R13129 a_n11737_n14973.n325 a_n11737_n14973.n324 4.5005
R13130 a_n11737_n14973.n118 a_n11737_n14973.n116 4.5005
R13131 a_n11737_n14973.n117 a_n11737_n14973.n323 4.5005
R13132 a_n11737_n14973.n322 a_n11737_n14973.n319 4.5005
R13133 a_n11737_n14973.n232 a_n11737_n14973.n224 4.5005
R13134 a_n11737_n14973.n112 a_n11737_n14973.n231 4.5005
R13135 a_n11737_n14973.n230 a_n11737_n14973.n111 4.5005
R13136 a_n11737_n14973.n229 a_n11737_n14973.n228 4.5005
R13137 a_n11737_n14973.n272 a_n11737_n14973.n271 4.5005
R13138 a_n11737_n14973.n270 a_n11737_n14973.n225 4.5005
R13139 a_n11737_n14973.n268 a_n11737_n14973.n267 4.5005
R13140 a_n11737_n14973.n266 a_n11737_n14973.n98 4.5005
R13141 a_n11737_n14973.n265 a_n11737_n14973.n100 4.5005
R13142 a_n11737_n14973.n99 a_n11737_n14973.n236 4.5005
R13143 a_n11737_n14973.n264 a_n11737_n14973.n263 4.5005
R13144 a_n11737_n14973.n252 a_n11737_n14973.n251 4.5005
R13145 a_n11737_n14973.n108 a_n11737_n14973.n253 4.5005
R13146 a_n11737_n14973.n254 a_n11737_n14973.n238 4.5005
R13147 a_n11737_n14973.n256 a_n11737_n14973.n255 4.5005
R13148 a_n11737_n14973.n257 a_n11737_n14973.n97 4.5005
R13149 a_n11737_n14973.n259 a_n11737_n14973.n258 4.5005
R13150 a_n11737_n14973.n260 a_n11737_n14973.n237 4.5005
R13151 a_n11737_n14973.n247 a_n11737_n14973.n246 4.5005
R13152 a_n11737_n14973.n245 a_n11737_n14973.n239 4.5005
R13153 a_n11737_n14973.n244 a_n11737_n14973.n243 4.5005
R13154 a_n11737_n14973.n242 a_n11737_n14973.n240 4.5005
R13155 a_n11737_n14973.n355 a_n11737_n14973.n141 4.5005
R13156 a_n11737_n14973.n134 a_n11737_n14973.n135 2.24296
R13157 a_n11737_n14973.n348 a_n11737_n14973.t10 3.83265
R13158 a_n11737_n14973.n344 a_n11737_n14973.n343 3.82765
R13159 a_n11737_n14973.n134 a_n11737_n14973.t16 3.82673
R13160 a_n11737_n14973.n354 a_n11737_n14973.n353 3.78255
R13161 a_n11737_n14973.n138 a_n11737_n14973.t26 3.76633
R13162 a_n11737_n14973.n359 a_n11737_n14973.n358 3.75068
R13163 a_n11737_n14973.n143 a_n11737_n14973.n142 3.75068
R13164 a_n11737_n14973.n356 a_n11737_n14973.t8 3.74975
R13165 a_n11737_n14973.n223 a_n11737_n14973.n145 3.37223
R13166 a_n11737_n14973.n113 a_n11737_n14973.n303 3.02216
R13167 a_n11737_n14973.n219 a_n11737_n14973.n218 2.89625
R13168 a_n11737_n14973.n18 a_n11737_n14973.n196 2.95081
R13169 a_n11737_n14973.n216 a_n11737_n14973.n161 2.88162
R13170 a_n11737_n14973.n194 a_n11737_n14973.n15 2.95081
R13171 a_n11737_n14973.n340 a_n11737_n14973.n339 2.76066
R13172 a_n11737_n14973.n339 a_n11737_n14973.n338 2.57313
R13173 a_n11737_n14973.n69 a_n11737_n14973.n83 2.00991
R13174 a_n11737_n14973.n274 a_n11737_n14973.n273 2.30989
R13175 a_n11737_n14973.n327 a_n11737_n14973.n146 2.30989
R13176 a_n11737_n14973.n303 a_n11737_n14973.n302 2.29659
R13177 a_n11737_n14973.n262 a_n11737_n14973.n261 2.2812
R13178 a_n11737_n14973.n357 a_n11737_n14973.n356 2.24389
R13179 a_n11737_n14973.n202 a_n11737_n14973.n172 2.23529
R13180 a_n11737_n14973.n184 a_n11737_n14973.n177 2.23529
R13181 a_n11737_n14973.n165 a_n11737_n14973.n163 2.23423
R13182 a_n11737_n14973.n157 a_n11737_n14973.n154 2.23423
R13183 a_n11737_n14973.n287 a_n11737_n14973.n275 2.18975
R13184 a_n11737_n14973.n326 a_n11737_n14973.n147 2.18975
R13185 a_n11737_n14973.n273 a_n11737_n14973.n224 2.16725
R13186 a_n11737_n14973.n252 a_n11737_n14973.n146 2.16725
R13187 a_n11737_n14973.n223 a_n11737_n14973.n222 2.11247
R13188 a_n11737_n14973.n188 a_n11737_n14973.n152 2.102
R13189 a_n11737_n14973.n46 a_n11737_n14973.n211 2.102
R13190 a_n11737_n14973.n352 a_n11737_n14973.n351 2.07395
R13191 a_n11737_n14973.n222 a_n11737_n14973.n152 2.07182
R13192 a_n11737_n14973.n212 a_n11737_n14973.n46 2.07182
R13193 a_n11737_n14973.n37 a_n11737_n14973.n66 2.13751
R13194 a_n11737_n14973.n213 a_n11737_n14973.n62 2.13751
R13195 a_n11737_n14973.n351 a_n11737_n14973.n340 1.90955
R13196 a_n11737_n14973.n333 a_n11737_n14973.n329 1.71486
R13197 a_n11737_n14973.n212 a_n11737_n14973.n145 1.50911
R13198 a_n11737_n14973.n222 a_n11737_n14973.n37 1.5005
R13199 a_n11737_n14973.n213 a_n11737_n14973.n212 1.5005
R13200 a_n11737_n14973.n275 a_n11737_n14973.n274 1.5005
R13201 a_n11737_n14973.n327 a_n11737_n14973.n326 1.5005
R13202 a_n11737_n14973.n333 a_n11737_n14973.n332 1.5005
R13203 a_n11737_n14973.n337 a_n11737_n14973.n336 1.5005
R13204 a_n11737_n14973.n351 a_n11737_n14973.n350 1.5005
R13205 a_n11737_n14973.n358 a_n11737_n14973.t13 1.4705
R13206 a_n11737_n14973.n358 a_n11737_n14973.t19 1.4705
R13207 a_n11737_n14973.n353 a_n11737_n14973.t21 1.4705
R13208 a_n11737_n14973.n353 a_n11737_n14973.t17 1.4705
R13209 a_n11737_n14973.n142 a_n11737_n14973.t24 1.4705
R13210 a_n11737_n14973.n142 a_n11737_n14973.t22 1.4705
R13211 a_n11737_n14973.n342 a_n11737_n14973.t20 1.4705
R13212 a_n11737_n14973.n342 a_n11737_n14973.t28 1.4705
R13213 a_n11737_n14973.n345 a_n11737_n14973.t11 1.4705
R13214 a_n11737_n14973.n345 a_n11737_n14973.t9 1.4705
R13215 a_n11737_n14973.n343 a_n11737_n14973.t27 1.4705
R13216 a_n11737_n14973.n343 a_n11737_n14973.t25 1.4705
R13217 a_n11737_n14973.n281 a_n11737_n14973.n280 1.39514
R13218 a_n11737_n14973.n274 a_n11737_n14973.n223 1.39023
R13219 a_n11737_n14973.n328 a_n11737_n14973.n327 1.39023
R13220 a_n11737_n14973.n144 a_n11737_n14973.n143 1.27228
R13221 a_n11737_n14973.n316 a_n11737_n14973.n315 1.26997
R13222 a_n11737_n14973.n289 a_n11737_n14973.n288 1.26997
R13223 a_n11737_n14973.n324 a_n11737_n14973.n318 1.24392
R13224 a_n11737_n14973.n292 a_n11737_n14973.n291 1.24392
R13225 a_n11737_n14973.n251 a_n11737_n14973.n250 1.24204
R13226 a_n11737_n14973.n233 a_n11737_n14973.n232 1.24204
R13227 a_n11737_n14973.n359 a_n11737_n14973.n357 1.20682
R13228 a_n11737_n14973.n248 a_n11737_n14973.n247 1.20414
R13229 a_n11737_n14973.n271 a_n11737_n14973.n235 1.20414
R13230 a_n11737_n14973.n322 a_n11737_n14973.n321 1.14132
R13231 a_n11737_n14973.n135 a_n11737_n14973.n354 1.20835
R13232 a_n11737_n14973.n229 a_n11737_n14973.n226 1.13598
R13233 a_n11737_n14973.n349 a_n11737_n14973.n344 1.13573
R13234 a_n11737_n14973.n335 a_n11737_n14973.n334 0.90675
R13235 a_n11737_n14973.n331 a_n11737_n14973.n330 0.90675
R13236 a_n11737_n14973.n344 a_n11737_n14973.n137 0.939226
R13237 a_n11737_n14973.n293 a_n11737_n14973.n275 0.752
R13238 a_n11737_n14973.n326 a_n11737_n14973.n325 0.752
R13239 a_n11737_n14973.n273 a_n11737_n14973.n272 0.71825
R13240 a_n11737_n14973.n246 a_n11737_n14973.n146 0.71825
R13241 a_n11737_n14973.n317 a_n11737_n14973.n316 0.663658
R13242 a_n11737_n14973.n318 a_n11737_n14973.n317 0.663658
R13243 a_n11737_n14973.n290 a_n11737_n14973.n289 0.663658
R13244 a_n11737_n14973.n291 a_n11737_n14973.n290 0.663658
R13245 a_n11737_n14973.n249 a_n11737_n14973.n248 0.655156
R13246 a_n11737_n14973.n250 a_n11737_n14973.n249 0.655156
R13247 a_n11737_n14973.n235 a_n11737_n14973.n234 0.655156
R13248 a_n11737_n14973.n234 a_n11737_n14973.n233 0.655156
R13249 a_n11737_n14973.n328 a_n11737_n14973.n145 0.603852
R13250 a_n11737_n14973.n354 a_n11737_n14973.n352 0.596867
R13251 a_n11737_n14973.n96 a_n11737_n14973.n95 0.313126
R13252 a_n11737_n14973.n280 a_n11737_n14973.n279 0.432797
R13253 a_n11737_n14973.n306 a_n11737_n14973.n114 0.394842
R13254 a_n11737_n14973.n301 a_n11737_n14973.n300 0.394842
R13255 a_n11737_n14973.n117 a_n11737_n14973.n319 0.381816
R13256 a_n11737_n14973.n296 a_n11737_n14973.n295 0.381816
R13257 a_n11737_n14973.n243 a_n11737_n14973.n242 0.379447
R13258 a_n11737_n14973.n260 a_n11737_n14973.n259 0.379447
R13259 a_n11737_n14973.n255 a_n11737_n14973.n254 0.379447
R13260 a_n11737_n14973.n268 a_n11737_n14973.n98 0.379447
R13261 a_n11737_n14973.n99 a_n11737_n14973.n264 0.379447
R13262 a_n11737_n14973.n228 a_n11737_n14973.n111 0.379447
R13263 a_n11737_n14973.n180 a_n11737_n14973.n52 0.44431
R13264 a_n11737_n14973.n79 a_n11737_n14973.n193 0.44431
R13265 a_n11737_n14973.n58 a_n11737_n14973.n173 0.44431
R13266 a_n11737_n14973.n1 a_n11737_n14973.n208 1.94004
R13267 a_n11737_n14973.n88 a_n11737_n14973.n105 0.44431
R13268 a_n11737_n14973.n94 a_n11737_n14973.n104 1.95665
R13269 a_n11737_n14973.n56 a_n11737_n14973.n179 0.44431
R13270 a_n11737_n14973.n80 a_n11737_n14973.n174 0.44431
R13271 a_n11737_n14973.n59 a_n11737_n14973.n197 0.44431
R13272 a_n11737_n14973.n299 a_n11737_n14973.n150 0.375125
R13273 a_n11737_n14973.n305 a_n11737_n14973.n304 0.375125
R13274 a_n11737_n14973.n192 a_n11737_n14973.n25 0.431935
R13275 a_n11737_n14973.n32 a_n11737_n14973.n207 0.431935
R13276 a_n11737_n14973.n73 a_n11737_n14973.n107 0.431935
R13277 a_n11737_n14973.n77 a_n11737_n14973.n106 0.431935
R13278 a_n11737_n14973.n29 a_n11737_n14973.n175 0.431935
R13279 a_n11737_n14973.n209 a_n11737_n14973.n33 0.431935
R13280 a_n11737_n14973.n297 a_n11737_n14973.n151 0.36275
R13281 a_n11737_n14973.n323 a_n11737_n14973.n322 0.36275
R13282 a_n11737_n14973.n185 a_n11737_n14973.n176 0.3605
R13283 a_n11737_n14973.n203 a_n11737_n14973.n171 0.3605
R13284 a_n11737_n14973.n158 a_n11737_n14973.n153 0.3605
R13285 a_n11737_n14973.n166 a_n11737_n14973.n164 0.3605
R13286 a_n11737_n14973.n38 a_n11737_n14973.n103 0.3605
R13287 a_n11737_n14973.n221 a_n11737_n14973.n72 0.429685
R13288 a_n11737_n14973.n220 a_n11737_n14973.n87 0.429685
R13289 a_n11737_n14973.n215 a_n11737_n14973.n214 0.3605
R13290 a_n11737_n14973.n170 a_n11737_n14973.n76 0.429685
R13291 a_n11737_n14973.n169 a_n11737_n14973.n94 1.93517
R13292 a_n11737_n14973.n230 a_n11737_n14973.n229 0.3605
R13293 a_n11737_n14973.n267 a_n11737_n14973.n266 0.3605
R13294 a_n11737_n14973.n263 a_n11737_n14973.n236 0.3605
R13295 a_n11737_n14973.n258 a_n11737_n14973.n237 0.3605
R13296 a_n11737_n14973.n256 a_n11737_n14973.n238 0.3605
R13297 a_n11737_n14973.n244 a_n11737_n14973.n240 0.3605
R13298 a_n11737_n14973.n352 a_n11737_n14973.n144 0.339591
R13299 a_n11737_n14973.n321 a_n11737_n14973.n320 0.335806
R13300 a_n11737_n14973.n227 a_n11737_n14973.n226 0.33475
R13301 a_n11737_n14973.n336 a_n11737_n14973.n335 0.320048
R13302 a_n11737_n14973.n332 a_n11737_n14973.n331 0.320048
R13303 a_n11737_n14973.n309 a_n11737_n14973.n148 0.302474
R13304 a_n11737_n14973.n284 a_n11737_n14973.n283 0.302474
R13305 a_n11737_n14973.n183 a_n11737_n14973.n182 0.287375
R13306 a_n11737_n14973.n199 a_n11737_n14973.n198 0.287375
R13307 a_n11737_n14973.n156 a_n11737_n14973.n155 0.287375
R13308 a_n11737_n14973.n162 a_n11737_n14973.n102 0.287375
R13309 a_n11737_n14973.n181 a_n11737_n14973.n178 0.287375
R13310 a_n11737_n14973.n47 a_n11737_n14973.n201 0.287375
R13311 a_n11737_n14973.n282 a_n11737_n14973.n277 0.287375
R13312 a_n11737_n14973.n311 a_n11737_n14973.n310 0.287375
R13313 a_n11737_n14973.n339 a_n11737_n14973.n337 0.212426
R13314 a_n11737_n14973.n158 a_n11737_n14973.n157 0.208888
R13315 a_n11737_n14973.n166 a_n11737_n14973.n163 0.208888
R13316 a_n11737_n14973.n185 a_n11737_n14973.n184 0.20887
R13317 a_n11737_n14973.n203 a_n11737_n14973.n202 0.20887
R13318 a_n11737_n14973.n357 a_n11737_n14973.n141 0.208385
R13319 a_n11737_n14973.n303 a_n11737_n14973.n150 0.208099
R13320 a_n11737_n14973.n262 a_n11737_n14973.n237 0.208099
R13321 a_n11737_n14973.n247 a_n11737_n14973.n239 0.147342
R13322 a_n11737_n14973.n259 a_n11737_n14973.n97 0.147342
R13323 a_n11737_n14973.n254 a_n11737_n14973.n108 0.147342
R13324 a_n11737_n14973.n271 a_n11737_n14973.n270 0.147342
R13325 a_n11737_n14973.n100 a_n11737_n14973.n98 0.147342
R13326 a_n11737_n14973.n112 a_n11737_n14973.n111 0.147342
R13327 a_n11737_n14973.n309 a_n11737_n14973.n308 0.147342
R13328 a_n11737_n14973.n313 a_n11737_n14973.n148 0.147342
R13329 a_n11737_n14973.n118 a_n11737_n14973.n117 0.147342
R13330 a_n11737_n14973.n283 a_n11737_n14973.n278 0.147342
R13331 a_n11737_n14973.n285 a_n11737_n14973.n284 0.147342
R13332 a_n11737_n14973.n295 a_n11737_n14973.n119 0.147342
R13333 a_n11737_n14973.n300 a_n11737_n14973.n101 0.147342
R13334 a_n11737_n14973.n139 a_n11737_n14973.n140 1.2061
R13335 a_n11737_n14973.n346 a_n11737_n14973.n139 0.230885
R13336 a_n11737_n14973.n346 a_n11737_n14973.n341 0.14
R13337 a_n11737_n14973.n136 a_n11737_n14973.n137 1.27228
R13338 a_n11737_n14973.t12 a_n11737_n14973.n136 6.50385
R13339 a_n11737_n14973.n182 a_n11737_n14973.n52 0.209185
R13340 a_n11737_n14973.n183 a_n11737_n14973.n44 0.209185
R13341 a_n11737_n14973.n184 a_n11737_n14973.n44 0.825446
R13342 a_n11737_n14973.n12 a_n11737_n14973.n176 0.209185
R13343 a_n11737_n14973.n7 a_n11737_n14973.n12 0.565419
R13344 a_n11737_n14973.n190 a_n11737_n14973.n7 0.834884
R13345 a_n11737_n14973.n191 a_n11737_n14973.n190 0.14
R13346 a_n11737_n14973.n192 a_n11737_n14973.n191 0.14
R13347 a_n11737_n14973.n193 a_n11737_n14973.n25 0.209185
R13348 a_n11737_n14973.n196 a_n11737_n14973.n79 0.209185
R13349 a_n11737_n14973.n18 a_n11737_n14973.n173 0.209185
R13350 a_n11737_n14973.n199 a_n11737_n14973.n58 0.209185
R13351 a_n11737_n14973.n198 a_n11737_n14973.n51 0.209185
R13352 a_n11737_n14973.n202 a_n11737_n14973.n51 0.825446
R13353 a_n11737_n14973.n14 a_n11737_n14973.n171 0.209185
R13354 a_n11737_n14973.n10 a_n11737_n14973.n14 0.565419
R13355 a_n11737_n14973.n205 a_n11737_n14973.n10 0.834884
R13356 a_n11737_n14973.n206 a_n11737_n14973.n205 0.14
R13357 a_n11737_n14973.n207 a_n11737_n14973.n206 0.14
R13358 a_n11737_n14973.n208 a_n11737_n14973.n32 0.209185
R13359 a_n11737_n14973.n155 a_n11737_n14973.n84 0.209185
R13360 a_n11737_n14973.n156 a_n11737_n14973.n41 0.209185
R13361 a_n11737_n14973.n157 a_n11737_n14973.n41 0.825427
R13362 a_n11737_n14973.n21 a_n11737_n14973.n153 0.209185
R13363 a_n11737_n14973.n160 a_n11737_n14973.n21 0.429685
R13364 a_n11737_n14973.n160 a_n11737_n14973.n129 0.208907
R13365 a_n11737_n14973.n67 a_n11737_n14973.n129 0.836657
R13366 a_n11737_n14973.n67 a_n11737_n14973.n107 0.209185
R13367 a_n11737_n14973.n73 a_n11737_n14973.n105 0.209185
R13368 a_n11737_n14973.n88 a_n11737_n14973.n161 0.209185
R13369 a_n11737_n14973.n216 a_n11737_n14973.n3 0.209185
R13370 a_n11737_n14973.n3 a_n11737_n14973.n92 0.513496
R13371 a_n11737_n14973.n92 a_n11737_n14973.n102 0.209185
R13372 a_n11737_n14973.n36 a_n11737_n14973.n162 0.209185
R13373 a_n11737_n14973.n36 a_n11737_n14973.n163 0.825427
R13374 a_n11737_n14973.n24 a_n11737_n14973.n164 0.209185
R13375 a_n11737_n14973.n168 a_n11737_n14973.n24 0.429685
R13376 a_n11737_n14973.n168 a_n11737_n14973.n126 0.208907
R13377 a_n11737_n14973.n63 a_n11737_n14973.n126 0.836657
R13378 a_n11737_n14973.n63 a_n11737_n14973.n106 0.209185
R13379 a_n11737_n14973.n77 a_n11737_n14973.n104 0.209185
R13380 a_n11737_n14973.n83 a_n11737_n14973.n103 0.209185
R13381 a_n11737_n14973.n39 a_n11737_n14973.n38 0.209137
R13382 a_n11737_n14973.n39 a_n11737_n14973.n37 0.886485
R13383 a_n11737_n14973.n221 a_n11737_n14973.n66 0.209113
R13384 a_n11737_n14973.n220 a_n11737_n14973.n72 0.209185
R13385 a_n11737_n14973.n219 a_n11737_n14973.n87 0.209185
R13386 a_n11737_n14973.n218 a_n11737_n14973.n4 0.209185
R13387 a_n11737_n14973.n91 a_n11737_n14973.n4 0.498871
R13388 a_n11737_n14973.n215 a_n11737_n14973.n91 0.209185
R13389 a_n11737_n14973.n214 a_n11737_n14973.n35 0.209137
R13390 a_n11737_n14973.n213 a_n11737_n14973.n35 0.886485
R13391 a_n11737_n14973.n170 a_n11737_n14973.n62 0.209113
R13392 a_n11737_n14973.n169 a_n11737_n14973.n76 0.209185
R13393 a_n11737_n14973.n56 a_n11737_n14973.n181 0.209185
R13394 a_n11737_n14973.n45 a_n11737_n14973.n178 0.209185
R13395 a_n11737_n14973.n152 a_n11737_n14973.n45 0.908935
R13396 a_n11737_n14973.n188 a_n11737_n14973.n187 0.14
R13397 a_n11737_n14973.n187 a_n11737_n14973.n175 0.14
R13398 a_n11737_n14973.n29 a_n11737_n14973.n174 0.209185
R13399 a_n11737_n14973.n194 a_n11737_n14973.n80 0.209185
R13400 a_n11737_n14973.n197 a_n11737_n14973.n15 0.209185
R13401 a_n11737_n14973.n201 a_n11737_n14973.n59 0.209185
R13402 a_n11737_n14973.n48 a_n11737_n14973.n47 0.209185
R13403 a_n11737_n14973.n48 a_n11737_n14973.n46 0.908935
R13404 a_n11737_n14973.n211 a_n11737_n14973.n130 0.14
R13405 a_n11737_n14973.n209 a_n11737_n14973.n130 0.14
R13406 a_n11737_n14973.n33 a_n11737_n14973.n0 1.54288
R13407 a_n11737_n14973.n282 a_n11737_n14973.n281 0.14
R13408 a_n11737_n14973.n286 a_n11737_n14973.n277 0.14
R13409 a_n11737_n14973.n287 a_n11737_n14973.n286 0.14
R13410 a_n11737_n14973.n294 a_n11737_n14973.n293 0.14
R13411 a_n11737_n14973.n294 a_n11737_n14973.n151 0.14
R13412 a_n11737_n14973.n298 a_n11737_n14973.n297 0.14
R13413 a_n11737_n14973.n299 a_n11737_n14973.n298 0.14
R13414 a_n11737_n14973.n304 a_n11737_n14973.n113 0.208168
R13415 a_n11737_n14973.n305 a_n11737_n14973.n149 0.14
R13416 a_n11737_n14973.n310 a_n11737_n14973.n149 0.14
R13417 a_n11737_n14973.n312 a_n11737_n14973.n311 0.14
R13418 a_n11737_n14973.n312 a_n11737_n14973.n147 0.14
R13419 a_n11737_n14973.n325 a_n11737_n14973.n116 0.14
R13420 a_n11737_n14973.n323 a_n11737_n14973.n116 0.14
R13421 a_n11737_n14973.n231 a_n11737_n14973.n230 0.14
R13422 a_n11737_n14973.n231 a_n11737_n14973.n224 0.14
R13423 a_n11737_n14973.n272 a_n11737_n14973.n225 0.14
R13424 a_n11737_n14973.n267 a_n11737_n14973.n225 0.14
R13425 a_n11737_n14973.n266 a_n11737_n14973.n265 0.14
R13426 a_n11737_n14973.n265 a_n11737_n14973.n236 0.14
R13427 a_n11737_n14973.n263 a_n11737_n14973.n110 0.208168
R13428 a_n11737_n14973.n110 a_n11737_n14973.n262 3.03679
R13429 a_n11737_n14973.n258 a_n11737_n14973.n257 0.14
R13430 a_n11737_n14973.n257 a_n11737_n14973.n256 0.14
R13431 a_n11737_n14973.n253 a_n11737_n14973.n238 0.14
R13432 a_n11737_n14973.n253 a_n11737_n14973.n252 0.14
R13433 a_n11737_n14973.n246 a_n11737_n14973.n245 0.14
R13434 a_n11737_n14973.n245 a_n11737_n14973.n244 0.14
R13435 a_n11737_n14973.n96 a_n11737_n14973.n240 1.12911
R13436 a_n11737_n14973.n141 a_n11737_n14973.n135 0.230894
R13437 a_n11737_n14973.n355 a_n11737_n14973.n134 0.138586
R13438 a_n11737_n14973.n347 a_n11737_n14973.n138 0.137318
R13439 a_n11737_n14973.n228 a_n11737_n14973.n227 0.128395
R13440 a_n11737_n14973.n320 a_n11737_n14973.n319 0.128395
R13441 a_n11737_n14973.n243 a_n11737_n14973.n241 0.118921
R13442 a_n11737_n14973.n261 a_n11737_n14973.n260 0.118921
R13443 a_n11737_n14973.n269 a_n11737_n14973.n268 0.118921
R13444 a_n11737_n14973.n315 a_n11737_n14973.n314 0.114184
R13445 a_n11737_n14973.n288 a_n11737_n14973.n276 0.114184
R13446 a_n11737_n14973.n307 a_n11737_n14973.n306 0.113
R13447 a_n11737_n14973.n348 a_n11737_n14973.n347 0.110782
R13448 a_n11737_n14973.n356 a_n11737_n14973.n355 0.109514
R13449 a_n11737_n14973.n13 a_n11737_n14973.n204 0.109179
R13450 a_n11737_n14973.n11 a_n11737_n14973.n186 0.109179
R13451 a_n11737_n14973.n57 a_n11737_n14973.n16 0.107155
R13452 a_n11737_n14973.n78 a_n11737_n14973.n27 0.107155
R13453 a_n11737_n14973.n55 a_n11737_n14973.n53 0.107155
R13454 a_n11737_n14973.n337 a_n11737_n14973.n333 0.105095
R13455 a_n11737_n14973.n131 a_n11737_n14973.n31 0.103632
R13456 a_n11737_n14973.n28 a_n11737_n14973.n26 0.103632
R13457 a_n11737_n14973.n302 a_n11737_n14973.n301 0.103526
R13458 a_n11737_n14973.n22 a_n11737_n14973.n167 0.102991
R13459 a_n11737_n14973.n124 a_n11737_n14973.n23 0.102991
R13460 a_n11737_n14973.n19 a_n11737_n14973.n159 0.102991
R13461 a_n11737_n14973.n127 a_n11737_n14973.n20 0.102991
R13462 a_n11737_n14973.n350 a_n11737_n14973.n349 0.0995
R13463 a_n11737_n14973.n75 a_n11737_n14973.n60 0.0933826
R13464 a_n11737_n14973.n71 a_n11737_n14973.n64 0.0933826
R13465 a_n11737_n14973.n93 a_n11737_n14973.n74 0.092742
R13466 a_n11737_n14973.n90 a_n11737_n14973.n2 0.092742
R13467 a_n11737_n14973.n86 a_n11737_n14973.n70 0.092742
R13468 a_n11737_n14973.n82 a_n11737_n14973.n68 0.092742
R13469 a_n11737_n14973.n200 a_n11737_n14973.n49 0.0821726
R13470 a_n11737_n14973.n42 a_n11737_n14973.n54 0.0821726
R13471 a_n11737_n14973.n120 a_n11737_n14973.n89 0.0821726
R13472 a_n11737_n14973.n121 a_n11737_n14973.n81 0.0821726
R13473 a_n11737_n14973.n128 a_n11737_n14973.n127 0.0427776
R13474 a_n11737_n14973.n125 a_n11737_n14973.n124 0.0427776
R13475 a_n11737_n14973.n350 a_n11737_n14973.n341 0.041
R13476 a_n11737_n14973.n132 a_n11737_n14973.n131 0.0402153
R13477 a_n11737_n14973.n26 a_n11737_n14973.n133 0.0402153
R13478 a_n11737_n14973.n53 a_n11737_n14973.n122 0.0402153
R13479 a_n11737_n14973.n189 a_n11737_n14973.n133 0.0402153
R13480 a_n11737_n14973.n210 a_n11737_n14973.n132 0.0402153
R13481 a_n11737_n14973.n308 a_n11737_n14973.n307 0.0348421
R13482 a_n11737_n14973.n279 a_n11737_n14973.n278 0.0348421
R13483 a_n11737_n14973.n204 a_n11737_n14973.n172 0.0344623
R13484 a_n11737_n14973.n186 a_n11737_n14973.n177 0.0344623
R13485 a_n11737_n14973.n314 a_n11737_n14973.n313 0.0336579
R13486 a_n11737_n14973.n285 a_n11737_n14973.n276 0.0336579
R13487 a_n11737_n14973.n167 a_n11737_n14973.n165 0.0325285
R13488 a_n11737_n14973.n159 a_n11737_n14973.n154 0.0325285
R13489 a_n11737_n14973.n241 a_n11737_n14973.n239 0.0289211
R13490 a_n11737_n14973.n270 a_n11737_n14973.n269 0.0289211
R13491 a_n11737_n14973.n242 a_n11737_n14973.n95 0.166289
R13492 a_n11737_n14973.n115 a_n11737_n14973.n114 0.156816
R13493 a_n11737_n14973.n264 a_n11737_n14973.n109 0.156816
R13494 a_n11737_n14973.n9 a_n11737_n14973.n8 0.154009
R13495 a_n11737_n14973.n6 a_n11737_n14973.n5 0.154009
R13496 a_n11737_n14973.n292 a_n11737_n14973.n119 0.147342
R13497 a_n11737_n14973.n324 a_n11737_n14973.n118 0.147342
R13498 a_n11737_n14973.n232 a_n11737_n14973.n112 0.147342
R13499 a_n11737_n14973.n251 a_n11737_n14973.n108 0.147342
R13500 a_n11737_n14973.n296 a_n11737_n14973.n101 0.147342
R13501 a_n11737_n14973.n100 a_n11737_n14973.n99 0.147342
R13502 a_n11737_n14973.n255 a_n11737_n14973.n97 0.147342
R13503 a_n11737_n14973.n90 a_n11737_n14973.n89 0.0943434
R13504 a_n11737_n14973.n82 a_n11737_n14973.n81 0.0943434
R13505 a_n11737_n14973.n75 a_n11737_n14973.n74 0.0901797
R13506 a_n11737_n14973.n71 a_n11737_n14973.n70 0.0901797
R13507 a_n11737_n14973.n8 a_n11737_n14973.n13 0.0847264
R13508 a_n11737_n14973.n5 a_n11737_n14973.n11 0.0847264
R13509 a_n11737_n14973.n86 a_n11737_n14973.n85 0.0799306
R13510 a_n11737_n14973.n195 a_n11737_n14973.n78 0.0799306
R13511 a_n11737_n14973.n65 a_n11737_n14973.n64 0.0799306
R13512 a_n11737_n14973.n61 a_n11737_n14973.n60 0.0799306
R13513 a_n11737_n14973.n200 a_n11737_n14973.n57 0.0799306
R13514 a_n11737_n14973.n55 a_n11737_n14973.n54 0.0799306
R13515 a_n11737_n14973.n50 a_n11737_n14973.n49 0.0799306
R13516 a_n11737_n14973.n43 a_n11737_n14973.n42 0.0799306
R13517 a_n11737_n14973.n121 a_n11737_n14973.n40 0.0799306
R13518 a_n11737_n14973.n120 a_n11737_n14973.n34 0.0799306
R13519 a_n11737_n14973.n31 a_n11737_n14973.n30 0.0799306
R13520 a_n11737_n14973.n28 a_n11737_n14973.n27 0.0799306
R13521 a_n11737_n14973.n23 a_n11737_n14973.n22 0.0799306
R13522 a_n11737_n14973.n20 a_n11737_n14973.n19 0.0799306
R13523 a_n11737_n14973.n17 a_n11737_n14973.n16 0.0799306
R13524 a_n11737_n14973.n217 a_n11737_n14973.n2 0.0799306
R13525 a_n11737_n14973.n1 a_n11737_n14973.t105 8.08727
C0 a_n1533_n16323# a_n1533_n16909# 0.008552f
C1 a_n965_n16909# a_n2101_n16909# 1.92e-19
C2 a_n965_n16909# a_n2631_n17634# 3.84e-20
C3 a_n2101_n16323# a_n2101_n16909# 0.008552f
C4 a_n1533_n16323# a_n965_n16909# 0.018349f
C5 a_n2101_n16323# a_n965_n16909# 1.92e-19
C6 a_n2101_n16323# a_n1533_n16323# 0.017228f
C7 a_n965_n15598# a_n965_n16909# 0.007268f
C8 a_n2631_n16323# a_n2631_n17634# 0.012404f
C9 a_n1533_n15598# a_n1533_n16323# 0.006281f
C10 a_n2631_n16323# a_n965_n16909# 3.84e-20
C11 AVDD IREF 0.25376p
C12 a_n1533_n15598# a_n965_n15598# 0.017228f
C13 a_n2101_n15598# a_n2101_n16323# 0.006281f
C14 a_n2631_n16323# a_n1533_n16323# 1.81e-19
C15 a_n2631_n16323# a_n2101_n16323# 0.017843f
C16 a_n2101_n15598# a_n1533_n15598# 0.017228f
C17 a_n2631_n16323# a_n965_n15598# 9.58e-21
C18 a_n1533_n17634# AVDD 0.04859f
C19 AVDD VN 70.0646f
C20 IREF VP 0.039954f
C21 a_n2631_n16323# a_n1533_n15598# 1.81e-19
C22 a_n2101_n17634# AVDD 0.030666f
C23 a_n2631_n16323# a_n2101_n15598# 0.017843f
C24 a_n1533_n16909# AVDD 0.016884f
C25 a_n2101_n16909# AVDD 0.016856f
C26 VP VN 55.8707f
C27 a_n2631_n17634# AVDD 0.378896f
C28 a_n965_n16909# AVDD 0.328969f
C29 a_n1533_n16323# AVDD 0.016884f
C30 a_n2101_n16323# AVDD 0.016856f
C31 a_n965_n15598# AVDD 0.165281f
C32 a_n1533_n15598# AVDD 0.030148f
C33 a_n2101_n15598# AVDD 0.030305f
C34 a_n2631_n16323# AVDD 0.378914f
C35 a_n6139_n20820# a_n6139_n21443# 0.007809f
C36 a_n6661_n21443# a_n6139_n21443# 0.017917f
C37 a_n6661_n21443# a_n6139_n20820# 0.017917f
C38 a_n5579_n20820# a_n6139_n20820# 0.017917f
C39 AVDD VP 63.8974f
C40 a_n5579_n20820# a_n6661_n21443# 2.78e-19
C41 a_n6139_n20267# a_n6139_n20820# 0.009337f
C42 a_n6139_n20267# a_n5579_n20820# 0.017917f
C43 a_n1533_n17634# IREF 0.001414f
C44 IREF VN 0.05459f
C45 AVDD VOUT 41.1792f
C46 a_n2101_n17634# IREF 0.001414f
C47 a_n2101_n17634# a_n1533_n17634# 0.017228f
C48 a_n2631_n17634# IREF 0.001629f
C49 a_n1533_n16909# a_n1533_n17634# 0.006281f
C50 a_n2101_n16909# a_n2101_n17634# 0.006281f
C51 a_n2631_n17634# a_n1533_n17634# 1.81e-19
C52 a_n2101_n16909# a_n1533_n16909# 0.017228f
C53 a_n2631_n17634# a_n2101_n17634# 0.017843f
C54 a_n2631_n17634# a_n1533_n16909# 1.81e-19
C55 a_n965_n16909# a_n1533_n16909# 0.018349f
C56 a_n2631_n17634# a_n2101_n16909# 0.017843f
C57 VOUT AVSS 13.120655f
C58 VN AVSS 18.261318f
C59 VP AVSS 18.257004f
C60 IREF AVSS 56.833004f
C61 AVDD AVSS 3.783745p
C62 a_n6139_n21443# AVSS 0.05176f
C63 a_n6139_n20820# AVSS 0.017025f
C64 a_n6661_n21443# AVSS 0.399052f
C65 a_n5579_n20820# AVSS 0.376201f
C66 a_n6139_n20267# AVSS 0.033958f
C67 a_n2631_n17634# AVSS 0.01042f
C68 a_n965_n16909# AVSS 0.010763f
C69 a_n965_n15598# AVSS 0.005065f
C70 a_n2631_n16323# AVSS 0.01042f
C71 a_n11737_n14973.n0 AVSS 0.053959f
C72 a_n11737_n14973.n1 AVSS 0.200819f
C73 a_n11737_n14973.n2 AVSS 0.168672f
C74 a_n11737_n14973.n3 AVSS 0.028681f
C75 a_n11737_n14973.n4 AVSS 0.028082f
C76 a_n11737_n14973.n5 AVSS 0.162298f
C77 a_n11737_n14973.n6 AVSS 0.194369f
C78 a_n11737_n14973.n7 AVSS 0.056804f
C79 a_n11737_n14973.n8 AVSS 0.162298f
C80 a_n11737_n14973.n9 AVSS 0.194369f
C81 a_n11737_n14973.n10 AVSS 0.056804f
C82 a_n11737_n14973.n11 AVSS 0.067733f
C83 a_n11737_n14973.n12 AVSS 0.031398f
C84 a_n11737_n14973.n13 AVSS 0.067733f
C85 a_n11737_n14973.n14 AVSS 0.031398f
C86 a_n11737_n14973.n15 AVSS 0.128388f
C87 a_n11737_n14973.n16 AVSS 0.073925f
C88 a_n11737_n14973.n17 AVSS 0.130496f
C89 a_n11737_n14973.n18 AVSS 0.128388f
C90 a_n11737_n14973.n19 AVSS 0.071823f
C91 a_n11737_n14973.n20 AVSS 0.168672f
C92 a_n11737_n14973.n21 AVSS 0.024786f
C93 a_n11737_n14973.n22 AVSS 0.071823f
C94 a_n11737_n14973.n23 AVSS 0.168672f
C95 a_n11737_n14973.n24 AVSS 0.024786f
C96 a_n11737_n14973.n25 AVSS 0.024881f
C97 a_n11737_n14973.n26 AVSS 0.072146f
C98 a_n11737_n14973.n27 AVSS 0.073925f
C99 a_n11737_n14973.n28 AVSS 0.168996f
C100 a_n11737_n14973.n29 AVSS 0.024881f
C101 a_n11737_n14973.n30 AVSS 0.073925f
C102 a_n11737_n14973.n31 AVSS 0.168996f
C103 a_n11737_n14973.n32 AVSS 0.024881f
C104 a_n11737_n14973.n33 AVSS 0.10043f
C105 a_n11737_n14973.n34 AVSS 0.132415f
C106 a_n11737_n14973.n35 AVSS 0.043743f
C107 a_n11737_n14973.n36 AVSS 0.041475f
C108 a_n11737_n14973.n37 AVSS 0.124071f
C109 a_n11737_n14973.n38 AVSS 0.024232f
C110 a_n11737_n14973.n39 AVSS 0.043743f
C111 a_n11737_n14973.n40 AVSS 0.132415f
C112 a_n11737_n14973.n41 AVSS 0.041475f
C113 a_n11737_n14973.n42 AVSS 0.061307f
C114 a_n11737_n14973.n43 AVSS 0.129499f
C115 a_n11737_n14973.n44 AVSS 0.041476f
C116 a_n11737_n14973.n45 AVSS 0.04465f
C117 a_n11737_n14973.n46 AVSS 0.390815f
C118 a_n11737_n14973.n47 AVSS 0.021241f
C119 a_n11737_n14973.n48 AVSS 0.04465f
C120 a_n11737_n14973.n49 AVSS 0.061307f
C121 a_n11737_n14973.n50 AVSS 0.129499f
C122 a_n11737_n14973.n51 AVSS 0.041476f
C123 a_n11737_n14973.n52 AVSS 0.0254f
C124 a_n11737_n14973.n53 AVSS 0.073925f
C125 a_n11737_n14973.n54 AVSS 0.061307f
C126 a_n11737_n14973.n55 AVSS 0.170772f
C127 a_n11737_n14973.n56 AVSS 0.0254f
C128 a_n11737_n14973.n57 AVSS 0.170772f
C129 a_n11737_n14973.n58 AVSS 0.0254f
C130 a_n11737_n14973.n59 AVSS 0.0254f
C131 a_n11737_n14973.n60 AVSS 0.071823f
C132 a_n11737_n14973.n61 AVSS 0.134664f
C133 a_n11737_n14973.n62 AVSS 0.095102f
C134 a_n11737_n14973.n63 AVSS 0.041933f
C135 a_n11737_n14973.n64 AVSS 0.071823f
C136 a_n11737_n14973.n65 AVSS 0.134664f
C137 a_n11737_n14973.n66 AVSS 0.095102f
C138 a_n11737_n14973.n67 AVSS 0.041933f
C139 a_n11737_n14973.n68 AVSS 0.162299f
C140 a_n11737_n14973.n69 AVSS 0.089278f
C141 a_n11737_n14973.n70 AVSS 0.071823f
C142 a_n11737_n14973.n71 AVSS 0.168996f
C143 a_n11737_n14973.n72 AVSS 0.024786f
C144 a_n11737_n14973.n73 AVSS 0.024881f
C145 a_n11737_n14973.n74 AVSS 0.071823f
C146 a_n11737_n14973.n75 AVSS 0.168996f
C147 a_n11737_n14973.n76 AVSS 0.024786f
C148 a_n11737_n14973.n77 AVSS 0.024881f
C149 a_n11737_n14973.n78 AVSS 0.170772f
C150 a_n11737_n14973.n79 AVSS 0.0254f
C151 a_n11737_n14973.n80 AVSS 0.0254f
C152 a_n11737_n14973.n81 AVSS 0.068585f
C153 a_n11737_n14973.n82 AVSS 0.170771f
C154 a_n11737_n14973.n83 AVSS 0.085765f
C155 a_n11737_n14973.n84 AVSS 0.088293f
C156 a_n11737_n14973.n85 AVSS 0.041503f
C157 a_n11737_n14973.n86 AVSS 0.170771f
C158 a_n11737_n14973.n87 AVSS 0.024786f
C159 a_n11737_n14973.n88 AVSS 0.0254f
C160 a_n11737_n14973.n89 AVSS 0.068585f
C161 a_n11737_n14973.n90 AVSS 0.170771f
C162 a_n11737_n14973.n91 AVSS 0.028082f
C163 a_n11737_n14973.n92 AVSS 0.028681f
C164 a_n11737_n14973.n93 AVSS 0.161789f
C165 a_n11737_n14973.n94 AVSS 0.089396f
C166 a_n11737_n14973.n95 AVSS 0.08438f
C167 a_n11737_n14973.n96 AVSS 0.137699f
C168 a_n11737_n14973.n97 AVSS 0.068283f
C169 a_n11737_n14973.n98 AVSS 0.019425f
C170 a_n11737_n14973.n99 AVSS 0.018725f
C171 a_n11737_n14973.n100 AVSS 0.068283f
C172 a_n11737_n14973.n101 AVSS 0.068283f
C173 a_n11737_n14973.n102 AVSS 0.021241f
C174 a_n11737_n14973.n103 AVSS 0.024234f
C175 a_n11737_n14973.n104 AVSS 0.08809f
C176 a_n11737_n14973.n105 AVSS 0.028114f
C177 a_n11737_n14973.n106 AVSS 0.02762f
C178 a_n11737_n14973.n107 AVSS 0.02762f
C179 a_n11737_n14973.n108 AVSS 0.067933f
C180 a_n11737_n14973.n109 AVSS 0.07948f
C181 a_n11737_n14973.n110 AVSS 0.132278f
C182 a_n11737_n14973.n111 AVSS 0.019425f
C183 a_n11737_n14973.n112 AVSS 0.067933f
C184 a_n11737_n14973.n113 AVSS 0.131604f
C185 a_n11737_n14973.n114 AVSS 0.019994f
C186 a_n11737_n14973.n115 AVSS 0.076933f
C187 a_n11737_n14973.n116 AVSS 0.011421f
C188 a_n11737_n14973.n117 AVSS 0.019513f
C189 a_n11737_n14973.n118 AVSS 0.067845f
C190 a_n11737_n14973.n119 AVSS 0.067845f
C191 a_n11737_n14973.n120 AVSS 0.064543f
C192 a_n11737_n14973.n121 AVSS 0.064543f
C193 a_n11737_n14973.n122 AVSS 0.098144f
C194 a_n11737_n14973.n123 AVSS 0.041813f
C195 a_n11737_n14973.n124 AVSS 0.071823f
C196 a_n11737_n14973.n125 AVSS 0.130873f
C197 a_n11737_n14973.n126 AVSS 0.042145f
C198 a_n11737_n14973.n127 AVSS 0.071823f
C199 a_n11737_n14973.n128 AVSS 0.130873f
C200 a_n11737_n14973.n129 AVSS 0.042145f
C201 a_n11737_n14973.n130 AVSS 0.011421f
C202 a_n11737_n14973.n131 AVSS 0.072146f
C203 a_n11737_n14973.n132 AVSS 0.09782f
C204 a_n11737_n14973.n133 AVSS 0.09782f
C205 a_n11737_n14973.n134 AVSS 0.08629f
C206 a_n11737_n14973.n135 AVSS 0.058565f
C207 a_n11737_n14973.n136 AVSS 0.257867f
C208 a_n11737_n14973.n137 AVSS 0.156445f
C209 a_n11737_n14973.n138 AVSS 0.083182f
C210 a_n11737_n14973.n139 AVSS 0.058467f
C211 a_n11737_n14973.n140 AVSS 0.253293f
C212 a_n11737_n14973.n141 AVSS 0.019764f
C213 a_n11737_n14973.t15 AVSS 0.100066f
C214 a_n11737_n14973.t24 AVSS 0.019342f
C215 a_n11737_n14973.t22 AVSS 0.019342f
C216 a_n11737_n14973.n142 AVSS 0.074133f
C217 a_n11737_n14973.n143 AVSS 0.255318f
C218 a_n11737_n14973.t18 AVSS 0.073923f
C219 a_n11737_n14973.n144 AVSS 0.129584f
C220 a_n11737_n14973.n145 AVSS 1.04628f
C221 a_n11737_n14973.n146 AVSS 0.457772f
C222 a_n11737_n14973.n147 AVSS 0.09533f
C223 a_n11737_n14973.n148 AVSS 0.016581f
C224 a_n11737_n14973.n149 AVSS 0.011421f
C225 a_n11737_n14973.n150 AVSS 0.024793f
C226 a_n11737_n14973.n151 AVSS 0.02054f
C227 a_n11737_n14973.t97 AVSS 0.160639f
C228 a_n11737_n14973.n152 AVSS 0.390815f
C229 a_n11737_n14973.n153 AVSS 0.024234f
C230 a_n11737_n14973.t101 AVSS 0.160639f
C231 a_n11737_n14973.n154 AVSS 0.133887f
C232 a_n11737_n14973.t58 AVSS 0.160639f
C233 a_n11737_n14973.t41 AVSS 0.160639f
C234 a_n11737_n14973.n155 AVSS 0.021241f
C235 a_n11737_n14973.n156 AVSS 0.021241f
C236 a_n11737_n14973.t66 AVSS 0.160639f
C237 a_n11737_n14973.n157 AVSS 0.041903f
C238 a_n11737_n14973.n158 AVSS 0.024223f
C239 a_n11737_n14973.n159 AVSS 0.06794f
C240 a_n11737_n14973.t86 AVSS 0.160639f
C241 a_n11737_n14973.n160 AVSS 0.02752f
C242 a_n11737_n14973.t102 AVSS 0.160639f
C243 a_n11737_n14973.t81 AVSS 0.160639f
C244 a_n11737_n14973.t53 AVSS 0.160639f
C245 a_n11737_n14973.n161 AVSS 0.127508f
C246 a_n11737_n14973.t82 AVSS 0.160639f
C247 a_n11737_n14973.t100 AVSS 0.160639f
C248 a_n11737_n14973.t80 AVSS 0.160639f
C249 a_n11737_n14973.n162 AVSS 0.021241f
C250 a_n11737_n14973.n163 AVSS 0.041903f
C251 a_n11737_n14973.t30 AVSS 0.160639f
C252 a_n11737_n14973.n164 AVSS 0.024234f
C253 a_n11737_n14973.t63 AVSS 0.160639f
C254 a_n11737_n14973.n165 AVSS 0.133887f
C255 a_n11737_n14973.n166 AVSS 0.024223f
C256 a_n11737_n14973.n167 AVSS 0.06794f
C257 a_n11737_n14973.t50 AVSS 0.160639f
C258 a_n11737_n14973.n168 AVSS 0.02752f
C259 a_n11737_n14973.t64 AVSS 0.160639f
C260 a_n11737_n14973.t73 AVSS 0.160639f
C261 a_n11737_n14973.t49 AVSS 0.160639f
C262 a_n11737_n14973.t74 AVSS 0.160639f
C263 a_n11737_n14973.n169 AVSS 0.090276f
C264 a_n11737_n14973.n170 AVSS 0.027528f
C265 a_n11737_n14973.n171 AVSS 0.024234f
C266 a_n11737_n14973.t45 AVSS 0.160639f
C267 a_n11737_n14973.n172 AVSS 0.129466f
C268 a_n11737_n14973.n173 AVSS 0.028114f
C269 a_n11737_n14973.t31 AVSS 0.160639f
C270 a_n11737_n14973.t44 AVSS 0.160639f
C271 a_n11737_n14973.n174 AVSS 0.028114f
C272 a_n11737_n14973.t84 AVSS 0.160639f
C273 a_n11737_n14973.n175 AVSS 0.023834f
C274 a_n11737_n14973.n176 AVSS 0.024234f
C275 a_n11737_n14973.t78 AVSS 0.160639f
C276 a_n11737_n14973.n177 AVSS 0.129466f
C277 a_n11737_n14973.t99 AVSS 0.160639f
C278 a_n11737_n14973.n178 AVSS 0.021241f
C279 a_n11737_n14973.t67 AVSS 0.160639f
C280 a_n11737_n14973.n179 AVSS 0.080208f
C281 a_n11737_n14973.t90 AVSS 0.160639f
C282 a_n11737_n14973.n180 AVSS 0.080199f
C283 a_n11737_n14973.n181 AVSS 0.021241f
C284 a_n11737_n14973.n182 AVSS 0.021241f
C285 a_n11737_n14973.n183 AVSS 0.021241f
C286 a_n11737_n14973.n184 AVSS 0.041903f
C287 a_n11737_n14973.n185 AVSS 0.024223f
C288 a_n11737_n14973.n186 AVSS 0.064072f
C289 a_n11737_n14973.t57 AVSS 0.160639f
C290 a_n11737_n14973.t79 AVSS 0.160639f
C291 a_n11737_n14973.t32 AVSS 0.160639f
C292 a_n11737_n14973.n187 AVSS 0.011421f
C293 a_n11737_n14973.n188 AVSS 0.091738f
C294 a_n11737_n14973.n189 AVSS 0.032676f
C295 a_n11737_n14973.n190 AVSS 0.040547f
C296 a_n11737_n14973.n191 AVSS 0.011421f
C297 a_n11737_n14973.n192 AVSS 0.023834f
C298 a_n11737_n14973.n193 AVSS 0.028114f
C299 a_n11737_n14973.t33 AVSS 0.160639f
C300 a_n11737_n14973.n194 AVSS 0.130339f
C301 a_n11737_n14973.n195 AVSS 0.033f
C302 a_n11737_n14973.n196 AVSS 0.130339f
C303 a_n11737_n14973.n197 AVSS 0.028114f
C304 a_n11737_n14973.n198 AVSS 0.021241f
C305 a_n11737_n14973.n199 AVSS 0.021241f
C306 a_n11737_n14973.n200 AVSS 0.061307f
C307 a_n11737_n14973.n201 AVSS 0.021241f
C308 a_n11737_n14973.t55 AVSS 0.160639f
C309 a_n11737_n14973.n202 AVSS 0.041903f
C310 a_n11737_n14973.n203 AVSS 0.024223f
C311 a_n11737_n14973.n204 AVSS 0.064072f
C312 a_n11737_n14973.t34 AVSS 0.160639f
C313 a_n11737_n14973.t47 AVSS 0.160639f
C314 a_n11737_n14973.n205 AVSS 0.040547f
C315 a_n11737_n14973.n206 AVSS 0.011421f
C316 a_n11737_n14973.n207 AVSS 0.023834f
C317 a_n11737_n14973.t75 AVSS 0.160639f
C318 a_n11737_n14973.n208 AVSS 0.087379f
C319 a_n11737_n14973.t105 AVSS 0.160965f
C320 a_n11737_n14973.n209 AVSS 0.023834f
C321 a_n11737_n14973.t104 AVSS 0.160639f
C322 a_n11737_n14973.n210 AVSS 0.032676f
C323 a_n11737_n14973.n211 AVSS 0.091738f
C324 a_n11737_n14973.n212 AVSS 1.67631f
C325 a_n11737_n14973.n213 AVSS 0.124071f
C326 a_n11737_n14973.n214 AVSS 0.024232f
C327 a_n11737_n14973.n215 AVSS 0.024234f
C328 a_n11737_n14973.n216 AVSS 0.12744f
C329 a_n11737_n14973.n217 AVSS 0.040394f
C330 a_n11737_n14973.n218 AVSS 0.128085f
C331 a_n11737_n14973.n219 AVSS 0.128038f
C332 a_n11737_n14973.n220 AVSS 0.02753f
C333 a_n11737_n14973.n221 AVSS 0.027528f
C334 a_n11737_n14973.n222 AVSS 1.78757f
C335 a_n11737_n14973.n223 AVSS 1.27422f
C336 a_n11737_n14973.n224 AVSS 0.094409f
C337 a_n11737_n14973.n225 AVSS 0.011421f
C338 a_n11737_n14973.t54 AVSS 0.164252f
C339 a_n11737_n14973.n226 AVSS 0.134251f
C340 a_n11737_n14973.t40 AVSS 0.160639f
C341 a_n11737_n14973.n227 AVSS 0.082128f
C342 a_n11737_n14973.n228 AVSS 0.018725f
C343 a_n11737_n14973.n229 AVSS 0.094248f
C344 a_n11737_n14973.n230 AVSS 0.020448f
C345 a_n11737_n14973.n231 AVSS 0.011421f
C346 a_n11737_n14973.t60 AVSS 0.160639f
C347 a_n11737_n14973.n232 AVSS 0.054743f
C348 a_n11737_n14973.t36 AVSS 0.160639f
C349 a_n11737_n14973.n233 AVSS 0.130911f
C350 a_n11737_n14973.t94 AVSS 0.160639f
C351 a_n11737_n14973.n234 AVSS 0.106378f
C352 a_n11737_n14973.t37 AVSS 0.160639f
C353 a_n11737_n14973.n235 AVSS 0.129549f
C354 a_n11737_n14973.n236 AVSS 0.020448f
C355 a_n11737_n14973.n237 AVSS 0.024194f
C356 a_n11737_n14973.n238 AVSS 0.020448f
C357 a_n11737_n14973.t70 AVSS 0.160639f
C358 a_n11737_n14973.t103 AVSS 0.160639f
C359 a_n11737_n14973.n239 AVSS 0.006475f
C360 a_n11737_n14973.n240 AVSS 0.098416f
C361 a_n11737_n14973.t68 AVSS 0.160639f
C362 a_n11737_n14973.n241 AVSS 0.062158f
C363 a_n11737_n14973.t42 AVSS 0.160639f
C364 a_n11737_n14973.t69 AVSS 0.164571f
C365 a_n11737_n14973.n242 AVSS 0.019425f
C366 a_n11737_n14973.n243 AVSS 0.018375f
C367 a_n11737_n14973.n244 AVSS 0.020448f
C368 a_n11737_n14973.n245 AVSS 0.011421f
C369 a_n11737_n14973.n246 AVSS 0.035093f
C370 a_n11737_n14973.n247 AVSS 0.053655f
C371 a_n11737_n14973.t85 AVSS 0.160639f
C372 a_n11737_n14973.n248 AVSS 0.129549f
C373 a_n11737_n14973.t59 AVSS 0.160639f
C374 a_n11737_n14973.n249 AVSS 0.106378f
C375 a_n11737_n14973.t83 AVSS 0.160639f
C376 a_n11737_n14973.n250 AVSS 0.130911f
C377 a_n11737_n14973.n251 AVSS 0.054743f
C378 a_n11737_n14973.n252 AVSS 0.094409f
C379 a_n11737_n14973.n253 AVSS 0.011421f
C380 a_n11737_n14973.n254 AVSS 0.019425f
C381 a_n11737_n14973.n255 AVSS 0.018725f
C382 a_n11737_n14973.n256 AVSS 0.020448f
C383 a_n11737_n14973.n257 AVSS 0.011421f
C384 a_n11737_n14973.n258 AVSS 0.020448f
C385 a_n11737_n14973.n259 AVSS 0.019425f
C386 a_n11737_n14973.n260 AVSS 0.018375f
C387 a_n11737_n14973.t91 AVSS 0.160639f
C388 a_n11737_n14973.n261 AVSS 0.077255f
C389 a_n11737_n14973.n262 AVSS 0.132403f
C390 a_n11737_n14973.t72 AVSS 0.160639f
C391 a_n11737_n14973.n263 AVSS 0.024197f
C392 a_n11737_n14973.n264 AVSS 0.019425f
C393 a_n11737_n14973.t46 AVSS 0.160639f
C394 a_n11737_n14973.n265 AVSS 0.011421f
C395 a_n11737_n14973.n266 AVSS 0.020448f
C396 a_n11737_n14973.n267 AVSS 0.020448f
C397 a_n11737_n14973.n268 AVSS 0.018375f
C398 a_n11737_n14973.t71 AVSS 0.160639f
C399 a_n11737_n14973.n269 AVSS 0.062158f
C400 a_n11737_n14973.n270 AVSS 0.006475f
C401 a_n11737_n14973.n271 AVSS 0.053655f
C402 a_n11737_n14973.n272 AVSS 0.035093f
C403 a_n11737_n14973.n273 AVSS 0.457772f
C404 a_n11737_n14973.n274 AVSS 1.65425f
C405 a_n11737_n14973.n275 AVSS 0.120383f
C406 a_n11737_n14973.t89 AVSS 0.160639f
C407 a_n11737_n14973.n276 AVSS 0.062158f
C408 a_n11737_n14973.n277 AVSS 0.017454f
C409 a_n11737_n14973.n278 AVSS 0.006694f
C410 a_n11737_n14973.t56 AVSS 0.160639f
C411 a_n11737_n14973.n279 AVSS 0.078951f
C412 a_n11737_n14973.t76 AVSS 0.163084f
C413 a_n11737_n14973.n280 AVSS 0.124527f
C414 a_n11737_n14973.n281 AVSS 0.086282f
C415 a_n11737_n14973.n282 AVSS 0.017454f
C416 a_n11737_n14973.n283 AVSS 0.016581f
C417 a_n11737_n14973.n284 AVSS 0.016581f
C418 a_n11737_n14973.n285 AVSS 0.00665f
C419 a_n11737_n14973.n286 AVSS 0.011421f
C420 a_n11737_n14973.n287 AVSS 0.09533f
C421 a_n11737_n14973.n288 AVSS 0.054798f
C422 a_n11737_n14973.t87 AVSS 0.160639f
C423 a_n11737_n14973.n289 AVSS 0.131086f
C424 a_n11737_n14973.t62 AVSS 0.160639f
C425 a_n11737_n14973.n290 AVSS 0.105733f
C426 a_n11737_n14973.t88 AVSS 0.160639f
C427 a_n11737_n14973.n291 AVSS 0.130211f
C428 a_n11737_n14973.n292 AVSS 0.054711f
C429 a_n11737_n14973.n293 AVSS 0.036474f
C430 a_n11737_n14973.n294 AVSS 0.011421f
C431 a_n11737_n14973.n295 AVSS 0.019513f
C432 a_n11737_n14973.t65 AVSS 0.160639f
C433 a_n11737_n14973.n296 AVSS 0.018813f
C434 a_n11737_n14973.n297 AVSS 0.02054f
C435 a_n11737_n14973.n298 AVSS 0.011421f
C436 a_n11737_n14973.n299 AVSS 0.021046f
C437 a_n11737_n14973.n300 AVSS 0.019994f
C438 a_n11737_n14973.n301 AVSS 0.018375f
C439 a_n11737_n14973.t98 AVSS 0.160639f
C440 a_n11737_n14973.n302 AVSS 0.078044f
C441 a_n11737_n14973.n303 AVSS 0.131932f
C442 a_n11737_n14973.t39 AVSS 0.160639f
C443 a_n11737_n14973.n304 AVSS 0.024796f
C444 a_n11737_n14973.n305 AVSS 0.021046f
C445 a_n11737_n14973.n306 AVSS 0.018725f
C446 a_n11737_n14973.t96 AVSS 0.160639f
C447 a_n11737_n14973.n307 AVSS 0.062158f
C448 a_n11737_n14973.n308 AVSS 0.006694f
C449 a_n11737_n14973.n309 AVSS 0.016581f
C450 a_n11737_n14973.n310 AVSS 0.017454f
C451 a_n11737_n14973.n311 AVSS 0.017454f
C452 a_n11737_n14973.n312 AVSS 0.011421f
C453 a_n11737_n14973.n313 AVSS 0.00665f
C454 a_n11737_n14973.t43 AVSS 0.160639f
C455 a_n11737_n14973.n314 AVSS 0.062158f
C456 a_n11737_n14973.n315 AVSS 0.054798f
C457 a_n11737_n14973.t51 AVSS 0.160639f
C458 a_n11737_n14973.n316 AVSS 0.131086f
C459 a_n11737_n14973.t38 AVSS 0.160639f
C460 a_n11737_n14973.n317 AVSS 0.105733f
C461 a_n11737_n14973.t52 AVSS 0.160639f
C462 a_n11737_n14973.n318 AVSS 0.130211f
C463 a_n11737_n14973.n319 AVSS 0.018813f
C464 a_n11737_n14973.t93 AVSS 0.164334f
C465 a_n11737_n14973.t61 AVSS 0.160639f
C466 a_n11737_n14973.n320 AVSS 0.082259f
C467 a_n11737_n14973.n321 AVSS 0.137456f
C468 a_n11737_n14973.n322 AVSS 0.097198f
C469 a_n11737_n14973.n323 AVSS 0.02054f
C470 a_n11737_n14973.t92 AVSS 0.160639f
C471 a_n11737_n14973.n324 AVSS 0.054711f
C472 a_n11737_n14973.n325 AVSS 0.036474f
C473 a_n11737_n14973.n326 AVSS 0.120383f
C474 a_n11737_n14973.n327 AVSS 1.65425f
C475 a_n11737_n14973.n328 AVSS 2.36877f
C476 a_n11737_n14973.t3 AVSS 0.102179f
C477 a_n11737_n14973.t7 AVSS 0.092168f
C478 a_n11737_n14973.n329 AVSS 0.362194f
C479 a_n11737_n14973.t35 AVSS 0.198966f
C480 a_n11737_n14973.t48 AVSS 0.191548f
C481 a_n11737_n14973.n330 AVSS 0.2601f
C482 a_n11737_n14973.t2 AVSS 0.19155f
C483 a_n11737_n14973.n331 AVSS 0.126637f
C484 a_n11737_n14973.t6 AVSS 0.1948f
C485 a_n11737_n14973.n332 AVSS 0.135748f
C486 a_n11737_n14973.n333 AVSS 0.340511f
C487 a_n11737_n14973.t4 AVSS 0.198966f
C488 a_n11737_n14973.t0 AVSS 0.191548f
C489 a_n11737_n14973.n334 AVSS 0.2601f
C490 a_n11737_n14973.t95 AVSS 0.19155f
C491 a_n11737_n14973.n335 AVSS 0.126637f
C492 a_n11737_n14973.t77 AVSS 0.1948f
C493 a_n11737_n14973.n336 AVSS 0.135748f
C494 a_n11737_n14973.n337 AVSS 0.177384f
C495 a_n11737_n14973.t5 AVSS 0.103194f
C496 a_n11737_n14973.t1 AVSS 0.080347f
C497 a_n11737_n14973.n338 AVSS 0.303945f
C498 a_n11737_n14973.n339 AVSS 0.805961f
C499 a_n11737_n14973.n340 AVSS 3.01817f
C500 a_n11737_n14973.n341 AVSS 0.007369f
C501 a_n11737_n14973.t14 AVSS 0.07429f
C502 a_n11737_n14973.t20 AVSS 0.019342f
C503 a_n11737_n14973.t28 AVSS 0.019342f
C504 a_n11737_n14973.n342 AVSS 0.074583f
C505 a_n11737_n14973.t12 AVSS 0.100858f
C506 a_n11737_n14973.t27 AVSS 0.019342f
C507 a_n11737_n14973.t25 AVSS 0.019342f
C508 a_n11737_n14973.n343 AVSS 0.076721f
C509 a_n11737_n14973.n344 AVSS 0.131391f
C510 a_n11737_n14973.t23 AVSS 0.100472f
C511 a_n11737_n14973.t11 AVSS 0.019342f
C512 a_n11737_n14973.t9 AVSS 0.019342f
C513 a_n11737_n14973.n345 AVSS 0.074583f
C514 a_n11737_n14973.t26 AVSS 0.048984f
C515 a_n11737_n14973.n346 AVSS 0.016006f
C516 a_n11737_n14973.n347 AVSS 0.007928f
C517 a_n11737_n14973.t10 AVSS 0.050146f
C518 a_n11737_n14973.n348 AVSS 0.086558f
C519 a_n11737_n14973.n349 AVSS 0.051204f
C520 a_n11737_n14973.n350 AVSS 0.005711f
C521 a_n11737_n14973.n351 AVSS 2.04334f
C522 a_n11737_n14973.n352 AVSS 0.348236f
C523 a_n11737_n14973.t21 AVSS 0.019342f
C524 a_n11737_n14973.t17 AVSS 0.019342f
C525 a_n11737_n14973.n353 AVSS 0.076147f
C526 a_n11737_n14973.n354 AVSS 0.119308f
C527 a_n11737_n14973.t16 AVSS 0.05004f
C528 a_n11737_n14973.n355 AVSS 0.007929f
C529 a_n11737_n14973.t8 AVSS 0.0487f
C530 a_n11737_n14973.n356 AVSS 0.081918f
C531 a_n11737_n14973.n357 AVSS 0.057502f
C532 a_n11737_n14973.t13 AVSS 0.019342f
C533 a_n11737_n14973.t19 AVSS 0.019342f
C534 a_n11737_n14973.n358 AVSS 0.074133f
C535 a_n11737_n14973.n359 AVSS 0.253716f
C536 a_n11737_n14973.t29 AVSS 0.100396f
C537 VOUT.t25 AVSS 0.087094f
C538 VOUT.t86 AVSS 0.087094f
C539 VOUT.n0 AVSS 0.191481f
C540 VOUT.n1 AVSS 0.114273f
C541 VOUT.n2 AVSS 0.76543f
C542 VOUT.n3 AVSS 0.051427f
C543 VOUT.t64 AVSS 0.260439f
C544 VOUT.n4 AVSS 0.40412f
C545 VOUT.n5 AVSS 0.051427f
C546 VOUT.t12 AVSS 0.087094f
C547 VOUT.t69 AVSS 0.087094f
C548 VOUT.n6 AVSS 0.257572f
C549 VOUT.n7 AVSS 0.311598f
C550 VOUT.t49 AVSS 0.680615f
C551 VOUT.n8 AVSS 1.67545f
C552 VOUT.n9 AVSS 0.114273f
C553 VOUT.n10 AVSS 0.306492f
C554 VOUT.n11 AVSS 3.82555f
C555 VOUT.n12 AVSS 3.76542f
C556 VOUT.t58 AVSS 0.087094f
C557 VOUT.t37 AVSS 0.087094f
C558 VOUT.n13 AVSS 0.837145f
C559 VOUT.t87 AVSS 0.391593f
C560 VOUT.n14 AVSS 2.24599f
C561 VOUT.t45 AVSS 0.087094f
C562 VOUT.t44 AVSS 0.087094f
C563 VOUT.n15 AVSS 0.837145f
C564 VOUT.t23 AVSS 0.391593f
C565 VOUT.n16 AVSS 2.24599f
C566 VOUT.n17 AVSS 2.33159f
C567 VOUT.t80 AVSS 0.229457f
C568 VOUT.t81 AVSS 0.244322f
C569 VOUT.n18 AVSS 0.927547f
C570 VOUT.t74 AVSS 0.087094f
C571 VOUT.t24 AVSS 0.087094f
C572 VOUT.n19 AVSS 0.221006f
C573 VOUT.t76 AVSS 0.087094f
C574 VOUT.t26 AVSS 0.087094f
C575 VOUT.n20 AVSS 0.238515f
C576 VOUT.n21 AVSS 0.60535f
C577 VOUT.n22 AVSS 0.504469f
C578 VOUT.t3 AVSS 0.087094f
C579 VOUT.t2 AVSS 0.087094f
C580 VOUT.n23 AVSS 0.40218f
C581 VOUT.n24 AVSS 1.97299f
C582 VOUT.t65 AVSS 0.391593f
C583 VOUT.n25 AVSS 1.83922f
C584 VOUT.n26 AVSS 5.67475f
C585 VOUT.n27 AVSS 0.239627f
C586 VOUT.t21 AVSS 0.229457f
C587 VOUT.t22 AVSS 0.244322f
C588 VOUT.n28 AVSS 0.773579f
C589 VOUT.n29 AVSS 0.596082f
C590 VOUT.t53 AVSS 0.229457f
C591 VOUT.t56 AVSS 0.244322f
C592 VOUT.n30 AVSS 0.770371f
C593 VOUT.n31 AVSS 0.705143f
C594 VOUT.t82 AVSS 0.087094f
C595 VOUT.t78 AVSS 0.087094f
C596 VOUT.n32 AVSS 0.221006f
C597 VOUT.t84 AVSS 0.087094f
C598 VOUT.t79 AVSS 0.087094f
C599 VOUT.n33 AVSS 0.238515f
C600 VOUT.n34 AVSS 0.60535f
C601 VOUT.n35 AVSS 0.47279f
C602 VOUT.t14 AVSS 0.229457f
C603 VOUT.t16 AVSS 0.244322f
C604 VOUT.n36 AVSS 0.78187f
C605 VOUT.n37 AVSS 0.717897f
C606 VOUT.t40 AVSS 0.229457f
C607 VOUT.t41 AVSS 0.244322f
C608 VOUT.n38 AVSS 0.78187f
C609 VOUT.n39 AVSS 0.717922f
C610 VOUT.t35 AVSS 0.087094f
C611 VOUT.t59 AVSS 0.087094f
C612 VOUT.n40 AVSS 0.221006f
C613 VOUT.t36 AVSS 0.087094f
C614 VOUT.t60 AVSS 0.087094f
C615 VOUT.n41 AVSS 0.238515f
C616 VOUT.n42 AVSS 0.60535f
C617 VOUT.n43 AVSS 0.336635f
C618 VOUT.t51 AVSS 0.229457f
C619 VOUT.t55 AVSS 0.244322f
C620 VOUT.n44 AVSS 0.92663f
C621 VOUT.t11 AVSS 0.087094f
C622 VOUT.t6 AVSS 0.087094f
C623 VOUT.n45 AVSS 0.221006f
C624 VOUT.t13 AVSS 0.087094f
C625 VOUT.t7 AVSS 0.087094f
C626 VOUT.n46 AVSS 0.238515f
C627 VOUT.n47 AVSS 0.60535f
C628 VOUT.n48 AVSS 0.639533f
C629 VOUT.t72 AVSS 0.229457f
C630 VOUT.t75 AVSS 0.244322f
C631 VOUT.n49 AVSS 0.770371f
C632 VOUT.n50 AVSS 0.705143f
C633 VOUT.t54 AVSS 0.229457f
C634 VOUT.t57 AVSS 0.244322f
C635 VOUT.n51 AVSS 0.773579f
C636 VOUT.n52 AVSS 0.596082f
C637 VOUT.n53 AVSS 0.239627f
C638 VOUT.n54 AVSS 5.20223f
C639 VOUT.n55 AVSS 0.051427f
C640 VOUT.n56 AVSS 0.051427f
C641 VOUT.n57 AVSS 0.76543f
C642 VOUT.t32 AVSS 0.087094f
C643 VOUT.t62 AVSS 0.087094f
C644 VOUT.n58 AVSS 0.257572f
C645 VOUT.n59 AVSS 0.311598f
C646 VOUT.n60 AVSS 0.114273f
C647 VOUT.n61 AVSS 0.210684f
C648 VOUT.n62 AVSS 0.210688f
C649 VOUT.t30 AVSS 0.260439f
C650 VOUT.n63 AVSS 0.40412f
C651 VOUT.n64 AVSS 0.114273f
C652 VOUT.n65 AVSS 1.34788f
C653 VOUT.n66 AVSS 0.051427f
C654 VOUT.t77 AVSS 0.087094f
C655 VOUT.t20 AVSS 0.087094f
C656 VOUT.n67 AVSS 0.257572f
C657 VOUT.n68 AVSS 0.311598f
C658 VOUT.t71 AVSS 0.680615f
C659 VOUT.n69 AVSS 1.67545f
C660 VOUT.n70 AVSS 0.114273f
C661 VOUT.n71 AVSS 0.306492f
C662 VOUT.n72 AVSS 1.60129f
C663 VOUT.n73 AVSS 3.30074f
C664 VOUT.n74 AVSS 3.19947f
C665 VOUT.n75 AVSS 1.65432f
C666 VOUT.t66 AVSS 0.087094f
C667 VOUT.t48 AVSS 0.087094f
C668 VOUT.n76 AVSS 0.40218f
C669 VOUT.n77 AVSS 1.97299f
C670 VOUT.t10 AVSS 0.391593f
C671 VOUT.n78 AVSS 1.29733f
C672 VOUT.n79 AVSS 3.53661f
C673 VOUT.t73 AVSS 0.229457f
C674 VOUT.t70 AVSS 0.244322f
C675 VOUT.n80 AVSS 0.927547f
C676 VOUT.t52 AVSS 0.087094f
C677 VOUT.t34 AVSS 0.087094f
C678 VOUT.n81 AVSS 0.221006f
C679 VOUT.t50 AVSS 0.087094f
C680 VOUT.t33 AVSS 0.087094f
C681 VOUT.n82 AVSS 0.238515f
C682 VOUT.n83 AVSS 0.60535f
C683 VOUT.n84 AVSS 0.504469f
C684 VOUT.t31 AVSS 0.229457f
C685 VOUT.t29 AVSS 0.244322f
C686 VOUT.n85 AVSS 0.92663f
C687 VOUT.t19 AVSS 0.087094f
C688 VOUT.t1 AVSS 0.087094f
C689 VOUT.n86 AVSS 0.221006f
C690 VOUT.t18 AVSS 0.087094f
C691 VOUT.t0 AVSS 0.087094f
C692 VOUT.n87 AVSS 0.238515f
C693 VOUT.n88 AVSS 0.60535f
C694 VOUT.n89 AVSS 0.639533f
C695 VOUT.t47 AVSS 0.229457f
C696 VOUT.t46 AVSS 0.244322f
C697 VOUT.n90 AVSS 0.770371f
C698 VOUT.n91 AVSS 0.705143f
C699 VOUT.t5 AVSS 0.229457f
C700 VOUT.t4 AVSS 0.244322f
C701 VOUT.n92 AVSS 0.773579f
C702 VOUT.n93 AVSS 0.596082f
C703 VOUT.n94 AVSS 0.239627f
C704 VOUT.t63 AVSS 0.087094f
C705 VOUT.t28 AVSS 0.087094f
C706 VOUT.n95 AVSS 0.221006f
C707 VOUT.t61 AVSS 0.087094f
C708 VOUT.t27 AVSS 0.087094f
C709 VOUT.n96 AVSS 0.238515f
C710 VOUT.n97 AVSS 0.60535f
C711 VOUT.n98 AVSS 0.336635f
C712 VOUT.t85 AVSS 0.229457f
C713 VOUT.t83 AVSS 0.244322f
C714 VOUT.n99 AVSS 0.78187f
C715 VOUT.n100 AVSS 0.717922f
C716 VOUT.t43 AVSS 0.229457f
C717 VOUT.t42 AVSS 0.244322f
C718 VOUT.n101 AVSS 0.78187f
C719 VOUT.n102 AVSS 0.717897f
C720 VOUT.t9 AVSS 0.087094f
C721 VOUT.t68 AVSS 0.087094f
C722 VOUT.n103 AVSS 0.221006f
C723 VOUT.t8 AVSS 0.087094f
C724 VOUT.t67 AVSS 0.087094f
C725 VOUT.n104 AVSS 0.238515f
C726 VOUT.n105 AVSS 0.60535f
C727 VOUT.n106 AVSS 0.47279f
C728 VOUT.t39 AVSS 0.229457f
C729 VOUT.t38 AVSS 0.244322f
C730 VOUT.n107 AVSS 0.770371f
C731 VOUT.n108 AVSS 0.705143f
C732 VOUT.t17 AVSS 0.229457f
C733 VOUT.t15 AVSS 0.244322f
C734 VOUT.n109 AVSS 0.773579f
C735 VOUT.n110 AVSS 0.596082f
C736 VOUT.n111 AVSS 0.239627f
C737 VOUT.n112 AVSS 3.82555f
C738 VOUT.n113 AVSS 7.49654f
C739 VOUT.n114 AVSS 0.051427f
C740 VOUT.t105 AVSS 0.082947f
C741 VOUT.t89 AVSS 0.082947f
C742 VOUT.n115 AVSS 0.239724f
C743 VOUT.n116 AVSS 0.321939f
C744 VOUT.t104 AVSS 0.632908f
C745 VOUT.n117 AVSS 1.54063f
C746 VOUT.n118 AVSS 0.114273f
C747 VOUT.n119 AVSS 1.32494f
C748 VOUT.t102 AVSS 0.082947f
C749 VOUT.t88 AVSS 0.082947f
C750 VOUT.n120 AVSS 0.206726f
C751 VOUT.t95 AVSS 0.082947f
C752 VOUT.t100 AVSS 0.082947f
C753 VOUT.n121 AVSS 0.222668f
C754 VOUT.n122 AVSS 0.74417f
C755 VOUT.t103 AVSS 0.082947f
C756 VOUT.t97 AVSS 0.082947f
C757 VOUT.n123 AVSS 0.206726f
C758 VOUT.t96 AVSS 0.082947f
C759 VOUT.t90 AVSS 0.082947f
C760 VOUT.n124 AVSS 0.222668f
C761 VOUT.n125 AVSS 0.905231f
C762 VOUT.t98 AVSS 0.227991f
C763 VOUT.t91 AVSS 0.241902f
C764 VOUT.n126 AVSS 0.743442f
C765 VOUT.n127 AVSS 1.03873f
C766 VOUT.t101 AVSS 0.227991f
C767 VOUT.t94 AVSS 0.241902f
C768 VOUT.n128 AVSS 0.746649f
C769 VOUT.n129 AVSS 0.601059f
C770 VOUT.n130 AVSS 0.570682f
C771 VOUT.n131 AVSS 6.16285f
C772 VOUT.t99 AVSS 0.082947f
C773 VOUT.t92 AVSS 0.082947f
C774 VOUT.n132 AVSS 0.745653f
C775 VOUT.t93 AVSS 0.381272f
C776 VOUT.n133 AVSS 2.59627f
C777 VOUT.n134 AVSS 4.30143f
C778 VOUT.n135 AVSS 7.46656f
C779 VOUT.n136 AVSS 5.91349f
C780 VOUT.n137 AVSS 1.60129f
C781 VOUT.n138 AVSS 1.34788f
C782 VOUT.n139 AVSS 0.114273f
C783 VOUT.n140 AVSS 0.210688f
C784 VOUT.n141 AVSS 0.210684f
C785 VOUT.n142 AVSS 0.051427f
C786 VOUT.n143 AVSS 0.115835f
C787 a_5396_9163.n0 AVSS 2.49493f
C788 a_5396_9163.n1 AVSS 2.1823f
C789 a_5396_9163.n2 AVSS 1.4092f
C790 a_5396_9163.n3 AVSS 2.49493f
C791 a_5396_9163.n4 AVSS 2.1823f
C792 a_5396_9163.n5 AVSS 1.4092f
C793 a_5396_9163.n6 AVSS 2.60308f
C794 a_5396_9163.n7 AVSS 1.84117f
C795 a_5396_9163.n8 AVSS 1.75569f
C796 a_5396_9163.n9 AVSS 2.60308f
C797 a_5396_9163.n10 AVSS 1.84117f
C798 a_5396_9163.n11 AVSS 1.33931f
C799 a_5396_9163.t73 AVSS 0.254253f
C800 a_5396_9163.t84 AVSS 0.270725f
C801 a_5396_9163.n12 AVSS 1.02677f
C802 a_5396_9163.t64 AVSS 0.096506f
C803 a_5396_9163.t44 AVSS 0.096506f
C804 a_5396_9163.n13 AVSS 0.244889f
C805 a_5396_9163.t43 AVSS 0.096506f
C806 a_5396_9163.t39 AVSS 0.096506f
C807 a_5396_9163.n14 AVSS 0.264291f
C808 a_5396_9163.n15 AVSS 0.670768f
C809 a_5396_9163.n16 AVSS 0.708645f
C810 a_5396_9163.t4 AVSS 0.254253f
C811 a_5396_9163.t14 AVSS 0.270725f
C812 a_5396_9163.n17 AVSS 0.853622f
C813 a_5396_9163.n18 AVSS 0.781345f
C814 a_5396_9163.t16 AVSS 0.096506f
C815 a_5396_9163.t68 AVSS 0.096506f
C816 a_5396_9163.n19 AVSS 0.244889f
C817 a_5396_9163.t65 AVSS 0.096506f
C818 a_5396_9163.t2 AVSS 0.096506f
C819 a_5396_9163.n20 AVSS 0.264291f
C820 a_5396_9163.n21 AVSS 0.670768f
C821 a_5396_9163.n22 AVSS 0.373014f
C822 a_5396_9163.n23 AVSS 3.54522f
C823 a_5396_9163.n24 AVSS 6.27658f
C824 a_5396_9163.n25 AVSS 6.288f
C825 a_5396_9163.t45 AVSS 0.096506f
C826 a_5396_9163.t11 AVSS 0.096506f
C827 a_5396_9163.n26 AVSS 0.449206f
C828 a_5396_9163.t82 AVSS 0.43646f
C829 a_5396_9163.t31 AVSS 0.096506f
C830 a_5396_9163.t1 AVSS 0.096506f
C831 a_5396_9163.n27 AVSS 0.449206f
C832 a_5396_9163.t71 AVSS 0.79093f
C833 a_5396_9163.t33 AVSS 0.433911f
C834 a_5396_9163.n28 AVSS 2.03798f
C835 a_5396_9163.t3 AVSS 0.096506f
C836 a_5396_9163.t72 AVSS 0.096506f
C837 a_5396_9163.n29 AVSS 0.445642f
C838 a_5396_9163.n30 AVSS 2.18621f
C839 a_5396_9163.t77 AVSS 0.096506f
C840 a_5396_9163.t60 AVSS 0.096506f
C841 a_5396_9163.n31 AVSS 0.927611f
C842 a_5396_9163.t19 AVSS 0.433911f
C843 a_5396_9163.n32 AVSS 2.4887f
C844 a_5396_9163.n33 AVSS 2.58355f
C845 a_5396_9163.t78 AVSS 0.254253f
C846 a_5396_9163.t86 AVSS 0.270725f
C847 a_5396_9163.n34 AVSS 1.02778f
C848 a_5396_9163.t62 AVSS 0.096506f
C849 a_5396_9163.t41 AVSS 0.096506f
C850 a_5396_9163.n35 AVSS 0.244889f
C851 a_5396_9163.t66 AVSS 0.096506f
C852 a_5396_9163.t48 AVSS 0.096506f
C853 a_5396_9163.n36 AVSS 0.264291f
C854 a_5396_9163.n37 AVSS 0.670768f
C855 a_5396_9163.n38 AVSS 0.558985f
C856 a_5396_9163.n39 AVSS 0.265523f
C857 a_5396_9163.t22 AVSS 0.254253f
C858 a_5396_9163.t28 AVSS 0.270725f
C859 a_5396_9163.n40 AVSS 0.857176f
C860 a_5396_9163.n41 AVSS 0.660498f
C861 a_5396_9163.t47 AVSS 0.254253f
C862 a_5396_9163.t51 AVSS 0.270725f
C863 a_5396_9163.n42 AVSS 0.853622f
C864 a_5396_9163.n43 AVSS 0.781345f
C865 a_5396_9163.t12 AVSS 0.096506f
C866 a_5396_9163.t76 AVSS 0.096506f
C867 a_5396_9163.n44 AVSS 0.244889f
C868 a_5396_9163.t23 AVSS 0.096506f
C869 a_5396_9163.t80 AVSS 0.096506f
C870 a_5396_9163.n45 AVSS 0.264291f
C871 a_5396_9163.n46 AVSS 0.670768f
C872 a_5396_9163.n47 AVSS 0.523883f
C873 a_5396_9163.t49 AVSS 0.254253f
C874 a_5396_9163.t54 AVSS 0.270725f
C875 a_5396_9163.n48 AVSS 0.866363f
C876 a_5396_9163.n49 AVSS 0.795477f
C877 a_5396_9163.t0 AVSS 0.254253f
C878 a_5396_9163.t5 AVSS 0.270725f
C879 a_5396_9163.n50 AVSS 0.866363f
C880 a_5396_9163.n51 AVSS 0.795504f
C881 a_5396_9163.t69 AVSS 0.096506f
C882 a_5396_9163.t34 AVSS 0.096506f
C883 a_5396_9163.n52 AVSS 0.244889f
C884 a_5396_9163.t74 AVSS 0.096506f
C885 a_5396_9163.t38 AVSS 0.096506f
C886 a_5396_9163.n53 AVSS 0.264291f
C887 a_5396_9163.n54 AVSS 0.670768f
C888 a_5396_9163.n55 AVSS 0.373014f
C889 a_5396_9163.t35 AVSS 0.254253f
C890 a_5396_9163.t42 AVSS 0.270725f
C891 a_5396_9163.n56 AVSS 1.02677f
C892 a_5396_9163.t26 AVSS 0.096506f
C893 a_5396_9163.t6 AVSS 0.096506f
C894 a_5396_9163.n57 AVSS 0.244889f
C895 a_5396_9163.t32 AVSS 0.096506f
C896 a_5396_9163.t9 AVSS 0.096506f
C897 a_5396_9163.n58 AVSS 0.264291f
C898 a_5396_9163.n59 AVSS 0.670768f
C899 a_5396_9163.n60 AVSS 0.708645f
C900 a_5396_9163.t55 AVSS 0.254253f
C901 a_5396_9163.t61 AVSS 0.270725f
C902 a_5396_9163.n61 AVSS 0.853622f
C903 a_5396_9163.n62 AVSS 0.781345f
C904 a_5396_9163.t10 AVSS 0.254253f
C905 a_5396_9163.t18 AVSS 0.270725f
C906 a_5396_9163.n63 AVSS 0.857176f
C907 a_5396_9163.n64 AVSS 0.660498f
C908 a_5396_9163.n65 AVSS 0.265523f
C909 a_5396_9163.n66 AVSS 5.76441f
C910 a_5396_9163.n67 AVSS 3.65744f
C911 a_5396_9163.n68 AVSS 1.8321f
C912 a_5396_9163.n69 AVSS 4.20978f
C913 a_5396_9163.t29 AVSS 0.096506f
C914 a_5396_9163.t7 AVSS 0.096506f
C915 a_5396_9163.n70 AVSS 0.927611f
C916 a_5396_9163.t57 AVSS 0.433911f
C917 a_5396_9163.n71 AVSS 2.4887f
C918 a_5396_9163.n72 AVSS 1.83309f
C919 a_5396_9163.t40 AVSS 0.096506f
C920 a_5396_9163.t20 AVSS 0.096506f
C921 a_5396_9163.n73 AVSS 0.445642f
C922 a_5396_9163.n74 AVSS 2.18621f
C923 a_5396_9163.t67 AVSS 0.433911f
C924 a_5396_9163.n75 AVSS 1.43753f
C925 a_5396_9163.n76 AVSS 3.91879f
C926 a_5396_9163.t30 AVSS 0.254253f
C927 a_5396_9163.t24 AVSS 0.270725f
C928 a_5396_9163.n77 AVSS 1.02778f
C929 a_5396_9163.t8 AVSS 0.096506f
C930 a_5396_9163.t75 AVSS 0.096506f
C931 a_5396_9163.n78 AVSS 0.244889f
C932 a_5396_9163.t15 AVSS 0.096506f
C933 a_5396_9163.t56 AVSS 0.096506f
C934 a_5396_9163.n79 AVSS 0.264291f
C935 a_5396_9163.n80 AVSS 0.670768f
C936 a_5396_9163.n81 AVSS 0.558985f
C937 a_5396_9163.t37 AVSS 0.254253f
C938 a_5396_9163.t70 AVSS 0.270725f
C939 a_5396_9163.n82 AVSS 0.866363f
C940 a_5396_9163.n83 AVSS 0.795504f
C941 a_5396_9163.t83 AVSS 0.254253f
C942 a_5396_9163.t46 AVSS 0.270725f
C943 a_5396_9163.n84 AVSS 0.866363f
C944 a_5396_9163.n85 AVSS 0.795477f
C945 a_5396_9163.t53 AVSS 0.096506f
C946 a_5396_9163.t27 AVSS 0.096506f
C947 a_5396_9163.n86 AVSS 0.244889f
C948 a_5396_9163.t25 AVSS 0.096506f
C949 a_5396_9163.t17 AVSS 0.096506f
C950 a_5396_9163.n87 AVSS 0.264291f
C951 a_5396_9163.n88 AVSS 0.670768f
C952 a_5396_9163.n89 AVSS 0.523883f
C953 a_5396_9163.t79 AVSS 0.254253f
C954 a_5396_9163.t85 AVSS 0.270725f
C955 a_5396_9163.n90 AVSS 0.853622f
C956 a_5396_9163.n91 AVSS 0.781345f
C957 a_5396_9163.t59 AVSS 0.254253f
C958 a_5396_9163.t52 AVSS 0.270725f
C959 a_5396_9163.n92 AVSS 0.857176f
C960 a_5396_9163.n93 AVSS 0.660498f
C961 a_5396_9163.n94 AVSS 0.265523f
C962 a_5396_9163.n95 AVSS 4.23896f
C963 a_5396_9163.n96 AVSS 3.72499f
C964 a_5396_9163.t168 AVSS 0.741107f
C965 a_5396_9163.t97 AVSS 0.096506f
C966 a_5396_9163.t169 AVSS 0.096506f
C967 a_5396_9163.n97 AVSS 0.385769f
C968 a_5396_9163.n98 AVSS 2.61131f
C969 a_5396_9163.n99 AVSS 4.08593f
C970 a_5396_9163.t163 AVSS 0.096506f
C971 a_5396_9163.t159 AVSS 0.096506f
C972 a_5396_9163.n100 AVSS 0.289434f
C973 a_5396_9163.t162 AVSS 0.096506f
C974 a_5396_9163.t155 AVSS 0.096506f
C975 a_5396_9163.n101 AVSS 0.224325f
C976 a_5396_9163.n102 AVSS 0.92886f
C977 a_5396_9163.t107 AVSS 0.096506f
C978 a_5396_9163.t125 AVSS 0.096506f
C979 a_5396_9163.n103 AVSS 0.289434f
C980 a_5396_9163.t106 AVSS 0.096506f
C981 a_5396_9163.t124 AVSS 0.096506f
C982 a_5396_9163.n104 AVSS 0.224325f
C983 a_5396_9163.n105 AVSS 0.66619f
C984 a_5396_9163.n106 AVSS 1.34217f
C985 a_5396_9163.t154 AVSS 0.096506f
C986 a_5396_9163.t149 AVSS 0.096506f
C987 a_5396_9163.n107 AVSS 0.289434f
C988 a_5396_9163.t153 AVSS 0.096506f
C989 a_5396_9163.t148 AVSS 0.096506f
C990 a_5396_9163.n108 AVSS 0.224325f
C991 a_5396_9163.n109 AVSS 0.66619f
C992 a_5396_9163.n110 AVSS 1.0395f
C993 a_5396_9163.t143 AVSS 0.096506f
C994 a_5396_9163.t93 AVSS 0.096506f
C995 a_5396_9163.n111 AVSS 0.289434f
C996 a_5396_9163.t157 AVSS 0.096506f
C997 a_5396_9163.t141 AVSS 0.096506f
C998 a_5396_9163.n112 AVSS 0.224325f
C999 a_5396_9163.n113 AVSS 0.66619f
C1000 a_5396_9163.n114 AVSS 0.2762f
C1001 a_5396_9163.t145 AVSS 0.381521f
C1002 a_5396_9163.t136 AVSS 0.096506f
C1003 a_5396_9163.t102 AVSS 0.096506f
C1004 a_5396_9163.n115 AVSS 0.384925f
C1005 a_5396_9163.t120 AVSS 0.381521f
C1006 a_5396_9163.t115 AVSS 0.096506f
C1007 a_5396_9163.t113 AVSS 0.096506f
C1008 a_5396_9163.n116 AVSS 0.883158f
C1009 a_5396_9163.n117 AVSS 2.61268f
C1010 a_5396_9163.n118 AVSS 5.69457f
C1011 a_5396_9163.n119 AVSS 0.811644f
C1012 a_5396_9163.t114 AVSS 0.096506f
C1013 a_5396_9163.t139 AVSS 0.096506f
C1014 a_5396_9163.n120 AVSS 0.289434f
C1015 a_5396_9163.t165 AVSS 0.096506f
C1016 a_5396_9163.t138 AVSS 0.096506f
C1017 a_5396_9163.n121 AVSS 0.224325f
C1018 a_5396_9163.n122 AVSS 0.66619f
C1019 a_5396_9163.n123 AVSS 1.02519f
C1020 a_5396_9163.t175 AVSS 0.096506f
C1021 a_5396_9163.t99 AVSS 0.096506f
C1022 a_5396_9163.n124 AVSS 0.289434f
C1023 a_5396_9163.t174 AVSS 0.096506f
C1024 a_5396_9163.t98 AVSS 0.096506f
C1025 a_5396_9163.n125 AVSS 0.224325f
C1026 a_5396_9163.n126 AVSS 0.66619f
C1027 a_5396_9163.n127 AVSS 1.03952f
C1028 a_5396_9163.t122 AVSS 0.096506f
C1029 a_5396_9163.t135 AVSS 0.096506f
C1030 a_5396_9163.n128 AVSS 0.289434f
C1031 a_5396_9163.t105 AVSS 0.096506f
C1032 a_5396_9163.t133 AVSS 0.096506f
C1033 a_5396_9163.n129 AVSS 0.224325f
C1034 a_5396_9163.n130 AVSS 0.66619f
C1035 a_5396_9163.n131 AVSS 1.0395f
C1036 a_5396_9163.t91 AVSS 0.096506f
C1037 a_5396_9163.t110 AVSS 0.096506f
C1038 a_5396_9163.n132 AVSS 0.289434f
C1039 a_5396_9163.t166 AVSS 0.096506f
C1040 a_5396_9163.t160 AVSS 0.096506f
C1041 a_5396_9163.n133 AVSS 0.224325f
C1042 a_5396_9163.n134 AVSS 0.66619f
C1043 a_5396_9163.n135 AVSS 0.578247f
C1044 a_5396_9163.n136 AVSS 6.48516f
C1045 a_5396_9163.t109 AVSS 0.741107f
C1046 a_5396_9163.t137 AVSS 0.096506f
C1047 a_5396_9163.t128 AVSS 0.096506f
C1048 a_5396_9163.n137 AVSS 0.385769f
C1049 a_5396_9163.n138 AVSS 2.61131f
C1050 a_5396_9163.n139 AVSS 1.83143f
C1051 a_5396_9163.t112 AVSS 0.382226f
C1052 a_5396_9163.n140 AVSS 1.82253f
C1053 a_5396_9163.t170 AVSS 0.096506f
C1054 a_5396_9163.t164 AVSS 0.096506f
C1055 a_5396_9163.n141 AVSS 0.385769f
C1056 a_5396_9163.n142 AVSS 1.40837f
C1057 a_5396_9163.n143 AVSS 4.68224f
C1058 a_5396_9163.n144 AVSS 4.05818f
C1059 a_5396_9163.t104 AVSS 0.381521f
C1060 a_5396_9163.t92 AVSS 0.096506f
C1061 a_5396_9163.t158 AVSS 0.096506f
C1062 a_5396_9163.n145 AVSS 0.384925f
C1063 a_5396_9163.t173 AVSS 0.381521f
C1064 a_5396_9163.t150 AVSS 0.096506f
C1065 a_5396_9163.t167 AVSS 0.096506f
C1066 a_5396_9163.n146 AVSS 0.883158f
C1067 a_5396_9163.n147 AVSS 1.83319f
C1068 a_5396_9163.n148 AVSS 3.66084f
C1069 a_5396_9163.t146 AVSS 0.096506f
C1070 a_5396_9163.t126 AVSS 0.096506f
C1071 a_5396_9163.n149 AVSS 0.289434f
C1072 a_5396_9163.t147 AVSS 0.096506f
C1073 a_5396_9163.t172 AVSS 0.096506f
C1074 a_5396_9163.n150 AVSS 0.224325f
C1075 a_5396_9163.n151 AVSS 0.66619f
C1076 a_5396_9163.n152 AVSS 0.578247f
C1077 a_5396_9163.t144 AVSS 0.096506f
C1078 a_5396_9163.t151 AVSS 0.096506f
C1079 a_5396_9163.n153 AVSS 0.289434f
C1080 a_5396_9163.t152 AVSS 0.096506f
C1081 a_5396_9163.t96 AVSS 0.096506f
C1082 a_5396_9163.n154 AVSS 0.224325f
C1083 a_5396_9163.n155 AVSS 0.66619f
C1084 a_5396_9163.n156 AVSS 1.0395f
C1085 a_5396_9163.t111 AVSS 0.096506f
C1086 a_5396_9163.t156 AVSS 0.096506f
C1087 a_5396_9163.n157 AVSS 0.289434f
C1088 a_5396_9163.t116 AVSS 0.096506f
C1089 a_5396_9163.t142 AVSS 0.096506f
C1090 a_5396_9163.n158 AVSS 0.224325f
C1091 a_5396_9163.n159 AVSS 0.66619f
C1092 a_5396_9163.n160 AVSS 1.03952f
C1093 a_5396_9163.t100 AVSS 0.096506f
C1094 a_5396_9163.t132 AVSS 0.096506f
C1095 a_5396_9163.n161 AVSS 0.289434f
C1096 a_5396_9163.t101 AVSS 0.096506f
C1097 a_5396_9163.t134 AVSS 0.096506f
C1098 a_5396_9163.n162 AVSS 0.224325f
C1099 a_5396_9163.n163 AVSS 0.66619f
C1100 a_5396_9163.n164 AVSS 1.02519f
C1101 a_5396_9163.t94 AVSS 0.096506f
C1102 a_5396_9163.t161 AVSS 0.096506f
C1103 a_5396_9163.n165 AVSS 0.289434f
C1104 a_5396_9163.t95 AVSS 0.096506f
C1105 a_5396_9163.t131 AVSS 0.096506f
C1106 a_5396_9163.n166 AVSS 0.224325f
C1107 a_5396_9163.n167 AVSS 0.92886f
C1108 a_5396_9163.t90 AVSS 0.096506f
C1109 a_5396_9163.t171 AVSS 0.096506f
C1110 a_5396_9163.n168 AVSS 0.289434f
C1111 a_5396_9163.t127 AVSS 0.096506f
C1112 a_5396_9163.t121 AVSS 0.096506f
C1113 a_5396_9163.n169 AVSS 0.224325f
C1114 a_5396_9163.n170 AVSS 0.66619f
C1115 a_5396_9163.n171 AVSS 1.34217f
C1116 a_5396_9163.t129 AVSS 0.096506f
C1117 a_5396_9163.t130 AVSS 0.096506f
C1118 a_5396_9163.n172 AVSS 0.289434f
C1119 a_5396_9163.t140 AVSS 0.096506f
C1120 a_5396_9163.t117 AVSS 0.096506f
C1121 a_5396_9163.n173 AVSS 0.224325f
C1122 a_5396_9163.n174 AVSS 0.66619f
C1123 a_5396_9163.n175 AVSS 1.0395f
C1124 a_5396_9163.t88 AVSS 0.096506f
C1125 a_5396_9163.t123 AVSS 0.096506f
C1126 a_5396_9163.n176 AVSS 0.289434f
C1127 a_5396_9163.t89 AVSS 0.096506f
C1128 a_5396_9163.t108 AVSS 0.096506f
C1129 a_5396_9163.n177 AVSS 0.224325f
C1130 a_5396_9163.n178 AVSS 0.66619f
C1131 a_5396_9163.n179 AVSS 0.2762f
C1132 a_5396_9163.n180 AVSS 0.811644f
C1133 a_5396_9163.n181 AVSS 3.69485f
C1134 a_5396_9163.n182 AVSS 4.40155f
C1135 a_5396_9163.n183 AVSS 1.83143f
C1136 a_5396_9163.t118 AVSS 0.382226f
C1137 a_5396_9163.n184 AVSS 1.82253f
C1138 a_5396_9163.t103 AVSS 0.096506f
C1139 a_5396_9163.t119 AVSS 0.096506f
C1140 a_5396_9163.n185 AVSS 0.385769f
C1141 a_5396_9163.n186 AVSS 1.40837f
C1142 a_5396_9163.n187 AVSS 5.45248f
C1143 a_5396_9163.n188 AVSS 6.21472f
C1144 a_5396_9163.n189 AVSS 4.99178f
C1145 a_5396_9163.t81 AVSS 0.096506f
C1146 a_5396_9163.t21 AVSS 0.096506f
C1147 a_5396_9163.n190 AVSS 0.449206f
C1148 a_5396_9163.t13 AVSS 0.43646f
C1149 a_5396_9163.t36 AVSS 0.096506f
C1150 a_5396_9163.t63 AVSS 0.096506f
C1151 a_5396_9163.n191 AVSS 0.449206f
C1152 a_5396_9163.t58 AVSS 0.79093f
C1153 a_5396_9163.n192 AVSS 1.8321f
C1154 a_5396_9163.n193 AVSS 4.91447f
C1155 a_5396_9163.n194 AVSS 4.23896f
C1156 a_5396_9163.n195 AVSS 0.265523f
C1157 a_5396_9163.n196 AVSS 0.660498f
C1158 a_5396_9163.t50 AVSS 0.254253f
C1159 a_5396_9163.n197 AVSS 0.857176f
C1160 a_5396_9163.t87 AVSS 0.270725f
C1161 a_n13990_n5465.n0 AVSS 1.90664f
C1162 a_n13990_n5465.n1 AVSS 1.66772f
C1163 a_n13990_n5465.n2 AVSS 1.07692f
C1164 a_n13990_n5465.n3 AVSS 1.90664f
C1165 a_n13990_n5465.n4 AVSS 1.66772f
C1166 a_n13990_n5465.n5 AVSS 1.07692f
C1167 a_n13990_n5465.n6 AVSS 2.07561f
C1168 a_n13990_n5465.n7 AVSS 1.81408f
C1169 a_n13990_n5465.n8 AVSS 1.44954f
C1170 a_n13990_n5465.n9 AVSS 1.55335f
C1171 a_n13990_n5465.t98 AVSS 0.194302f
C1172 a_n13990_n5465.t99 AVSS 0.20689f
C1173 a_n13990_n5465.n10 AVSS 0.784662f
C1174 a_n13990_n5465.t27 AVSS 0.073751f
C1175 a_n13990_n5465.t74 AVSS 0.073751f
C1176 a_n13990_n5465.n11 AVSS 0.187146f
C1177 a_n13990_n5465.t29 AVSS 0.073751f
C1178 a_n13990_n5465.t75 AVSS 0.073751f
C1179 a_n13990_n5465.n12 AVSS 0.201973f
C1180 a_n13990_n5465.n13 AVSS 0.512605f
C1181 a_n13990_n5465.n14 AVSS 0.541551f
C1182 a_n13990_n5465.t101 AVSS 0.073751f
C1183 a_n13990_n5465.t81 AVSS 0.073751f
C1184 a_n13990_n5465.n15 AVSS 0.187146f
C1185 a_n13990_n5465.t105 AVSS 0.073751f
C1186 a_n13990_n5465.t82 AVSS 0.073751f
C1187 a_n13990_n5465.n16 AVSS 0.201973f
C1188 a_n13990_n5465.n17 AVSS 0.512605f
C1189 a_n13990_n5465.n18 AVSS 0.28506f
C1190 a_n13990_n5465.t32 AVSS 0.073751f
C1191 a_n13990_n5465.t94 AVSS 0.073751f
C1192 a_n13990_n5465.n19 AVSS 0.708887f
C1193 a_n13990_n5465.t93 AVSS 0.331597f
C1194 a_n13990_n5465.n20 AVSS 1.90188f
C1195 a_n13990_n5465.n21 AVSS 1.97437f
C1196 a_n13990_n5465.n22 AVSS 2.70928f
C1197 a_n13990_n5465.t70 AVSS 0.073751f
C1198 a_n13990_n5465.t43 AVSS 0.073751f
C1199 a_n13990_n5465.n23 AVSS 0.340562f
C1200 a_n13990_n5465.n24 AVSS 1.67071f
C1201 a_n13990_n5465.t61 AVSS 0.331597f
C1202 a_n13990_n5465.n25 AVSS 1.55743f
C1203 a_n13990_n5465.t52 AVSS 0.194302f
C1204 a_n13990_n5465.t53 AVSS 0.20689f
C1205 a_n13990_n5465.n26 AVSS 0.785438f
C1206 a_n13990_n5465.t42 AVSS 0.073751f
C1207 a_n13990_n5465.t34 AVSS 0.073751f
C1208 a_n13990_n5465.n27 AVSS 0.187146f
C1209 a_n13990_n5465.t44 AVSS 0.073751f
C1210 a_n13990_n5465.t35 AVSS 0.073751f
C1211 a_n13990_n5465.n28 AVSS 0.201973f
C1212 a_n13990_n5465.n29 AVSS 0.512605f
C1213 a_n13990_n5465.n30 AVSS 0.42718f
C1214 a_n13990_n5465.t40 AVSS 0.194302f
C1215 a_n13990_n5465.t41 AVSS 0.20689f
C1216 a_n13990_n5465.n31 AVSS 0.662081f
C1217 a_n13990_n5465.n32 AVSS 0.607929f
C1218 a_n13990_n5465.t46 AVSS 0.194302f
C1219 a_n13990_n5465.t49 AVSS 0.20689f
C1220 a_n13990_n5465.n33 AVSS 0.662081f
C1221 a_n13990_n5465.n34 AVSS 0.607909f
C1222 a_n13990_n5465.t83 AVSS 0.073751f
C1223 a_n13990_n5465.t37 AVSS 0.073751f
C1224 a_n13990_n5465.n35 AVSS 0.187146f
C1225 a_n13990_n5465.t85 AVSS 0.073751f
C1226 a_n13990_n5465.t39 AVSS 0.073751f
C1227 a_n13990_n5465.n36 AVSS 0.201973f
C1228 a_n13990_n5465.n37 AVSS 0.512605f
C1229 a_n13990_n5465.n38 AVSS 0.400355f
C1230 a_n13990_n5465.t78 AVSS 0.194302f
C1231 a_n13990_n5465.t79 AVSS 0.20689f
C1232 a_n13990_n5465.n39 AVSS 0.652343f
C1233 a_n13990_n5465.n40 AVSS 0.597109f
C1234 a_n13990_n5465.t91 AVSS 0.194302f
C1235 a_n13990_n5465.t92 AVSS 0.20689f
C1236 a_n13990_n5465.n41 AVSS 0.655059f
C1237 a_n13990_n5465.n42 AVSS 0.504757f
C1238 a_n13990_n5465.n43 AVSS 0.202914f
C1239 a_n13990_n5465.n44 AVSS 4.80533f
C1240 a_n13990_n5465.n45 AVSS 4.37207f
C1241 a_n13990_n5465.t38 AVSS 0.194302f
C1242 a_n13990_n5465.t36 AVSS 0.20689f
C1243 a_n13990_n5465.n46 AVSS 0.785438f
C1244 a_n13990_n5465.t90 AVSS 0.073751f
C1245 a_n13990_n5465.t65 AVSS 0.073751f
C1246 a_n13990_n5465.n47 AVSS 0.187146f
C1247 a_n13990_n5465.t89 AVSS 0.073751f
C1248 a_n13990_n5465.t63 AVSS 0.073751f
C1249 a_n13990_n5465.n48 AVSS 0.201973f
C1250 a_n13990_n5465.n49 AVSS 0.512605f
C1251 a_n13990_n5465.n50 AVSS 0.42718f
C1252 a_n13990_n5465.t103 AVSS 0.194302f
C1253 a_n13990_n5465.t100 AVSS 0.20689f
C1254 a_n13990_n5465.n51 AVSS 0.784662f
C1255 a_n13990_n5465.t51 AVSS 0.073751f
C1256 a_n13990_n5465.t107 AVSS 0.073751f
C1257 a_n13990_n5465.n52 AVSS 0.187146f
C1258 a_n13990_n5465.t50 AVSS 0.073751f
C1259 a_n13990_n5465.t106 AVSS 0.073751f
C1260 a_n13990_n5465.n53 AVSS 0.201973f
C1261 a_n13990_n5465.n54 AVSS 0.512605f
C1262 a_n13990_n5465.n55 AVSS 0.541551f
C1263 a_n13990_n5465.t25 AVSS 0.194302f
C1264 a_n13990_n5465.t111 AVSS 0.20689f
C1265 a_n13990_n5465.n56 AVSS 0.652343f
C1266 a_n13990_n5465.n57 AVSS 0.597109f
C1267 a_n13990_n5465.t86 AVSS 0.194302f
C1268 a_n13990_n5465.t84 AVSS 0.20689f
C1269 a_n13990_n5465.n58 AVSS 0.655059f
C1270 a_n13990_n5465.n59 AVSS 0.504757f
C1271 a_n13990_n5465.n60 AVSS 4.24693f
C1272 a_n13990_n5465.t119 AVSS 0.070239f
C1273 a_n13990_n5465.t17 AVSS 0.070239f
C1274 a_n13990_n5465.n61 AVSS 0.320902f
C1275 a_n13990_n5465.t120 AVSS 0.561285f
C1276 a_n13990_n5465.n62 AVSS 1.9181f
C1277 a_n13990_n5465.t141 AVSS 0.070239f
C1278 a_n13990_n5465.t22 AVSS 0.070239f
C1279 a_n13990_n5465.n63 AVSS 0.175054f
C1280 a_n13990_n5465.t139 AVSS 0.070239f
C1281 a_n13990_n5465.t12 AVSS 0.070239f
C1282 a_n13990_n5465.n64 AVSS 0.188553f
C1283 a_n13990_n5465.n65 AVSS 0.630156f
C1284 a_n13990_n5465.t116 AVSS 0.070239f
C1285 a_n13990_n5465.t140 AVSS 0.070239f
C1286 a_n13990_n5465.n66 AVSS 0.320902f
C1287 a_n13990_n5465.t117 AVSS 0.324757f
C1288 a_n13990_n5465.n67 AVSS 5.25784f
C1289 a_n13990_n5465.n68 AVSS 0.483248f
C1290 a_n13990_n5465.t11 AVSS 0.193061f
C1291 a_n13990_n5465.t0 AVSS 0.204841f
C1292 a_n13990_n5465.n69 AVSS 0.632256f
C1293 a_n13990_n5465.n70 AVSS 0.508971f
C1294 a_n13990_n5465.t8 AVSS 0.193061f
C1295 a_n13990_n5465.t15 AVSS 0.204841f
C1296 a_n13990_n5465.n71 AVSS 0.62954f
C1297 a_n13990_n5465.n72 AVSS 0.598514f
C1298 a_n13990_n5465.t3 AVSS 0.070239f
C1299 a_n13990_n5465.t9 AVSS 0.070239f
C1300 a_n13990_n5465.n73 AVSS 0.175054f
C1301 a_n13990_n5465.t1 AVSS 0.070239f
C1302 a_n13990_n5465.t16 AVSS 0.070239f
C1303 a_n13990_n5465.n74 AVSS 0.188553f
C1304 a_n13990_n5465.n75 AVSS 0.52607f
C1305 a_n13990_n5465.n76 AVSS 0.79473f
C1306 a_n13990_n5465.t113 AVSS 0.070239f
C1307 a_n13990_n5465.t7 AVSS 0.070239f
C1308 a_n13990_n5465.n77 AVSS 0.175054f
C1309 a_n13990_n5465.t118 AVSS 0.070239f
C1310 a_n13990_n5465.t24 AVSS 0.070239f
C1311 a_n13990_n5465.n78 AVSS 0.188553f
C1312 a_n13990_n5465.n79 AVSS 0.52607f
C1313 a_n13990_n5465.n80 AVSS 0.679337f
C1314 a_n13990_n5465.t13 AVSS 0.070239f
C1315 a_n13990_n5465.t19 AVSS 0.070239f
C1316 a_n13990_n5465.n81 AVSS 0.175054f
C1317 a_n13990_n5465.t20 AVSS 0.070239f
C1318 a_n13990_n5465.t6 AVSS 0.070239f
C1319 a_n13990_n5465.n82 AVSS 0.188553f
C1320 a_n13990_n5465.n83 AVSS 0.766542f
C1321 a_n13990_n5465.t18 AVSS 0.193061f
C1322 a_n13990_n5465.t5 AVSS 0.204841f
C1323 a_n13990_n5465.n84 AVSS 0.62954f
C1324 a_n13990_n5465.n85 AVSS 0.879586f
C1325 a_n13990_n5465.t23 AVSS 0.193061f
C1326 a_n13990_n5465.t4 AVSS 0.204841f
C1327 a_n13990_n5465.n86 AVSS 0.632256f
C1328 a_n13990_n5465.n87 AVSS 0.508971f
C1329 a_n13990_n5465.n88 AVSS 0.20023f
C1330 a_n13990_n5465.n89 AVSS 4.63877f
C1331 a_n13990_n5465.t114 AVSS 0.322858f
C1332 a_n13990_n5465.n90 AVSS 1.05136f
C1333 a_n13990_n5465.t2 AVSS 0.070239f
C1334 a_n13990_n5465.t115 AVSS 0.070239f
C1335 a_n13990_n5465.n91 AVSS 0.318412f
C1336 a_n13990_n5465.n92 AVSS 1.47152f
C1337 a_n13990_n5465.t14 AVSS 0.070239f
C1338 a_n13990_n5465.t10 AVSS 0.070239f
C1339 a_n13990_n5465.n93 AVSS 0.631412f
C1340 a_n13990_n5465.t21 AVSS 0.322858f
C1341 a_n13990_n5465.n94 AVSS 1.82196f
C1342 a_n13990_n5465.n95 AVSS 1.19295f
C1343 a_n13990_n5465.n96 AVSS 4.80062f
C1344 a_n13990_n5465.n97 AVSS 5.18898f
C1345 a_n13990_n5465.t126 AVSS 0.284312f
C1346 a_n13990_n5465.t124 AVSS 0.070239f
C1347 a_n13990_n5465.t125 AVSS 0.070239f
C1348 a_n13990_n5465.n98 AVSS 0.595322f
C1349 a_n13990_n5465.n99 AVSS 3.49889f
C1350 a_n13990_n5465.t132 AVSS 0.219819f
C1351 a_n13990_n5465.t133 AVSS 0.180853f
C1352 a_n13990_n5465.n100 AVSS 0.786008f
C1353 a_n13990_n5465.t121 AVSS 0.070239f
C1354 a_n13990_n5465.t130 AVSS 0.070239f
C1355 a_n13990_n5465.n101 AVSS 0.205803f
C1356 a_n13990_n5465.t134 AVSS 0.070239f
C1357 a_n13990_n5465.t131 AVSS 0.070239f
C1358 a_n13990_n5465.n102 AVSS 0.161282f
C1359 a_n13990_n5465.n103 AVSS 0.522594f
C1360 a_n13990_n5465.n104 AVSS 0.967708f
C1361 a_n13990_n5465.t123 AVSS 0.070239f
C1362 a_n13990_n5465.t136 AVSS 0.070239f
C1363 a_n13990_n5465.n105 AVSS 0.205803f
C1364 a_n13990_n5465.t135 AVSS 0.070239f
C1365 a_n13990_n5465.t127 AVSS 0.070239f
C1366 a_n13990_n5465.n106 AVSS 0.161282f
C1367 a_n13990_n5465.n107 AVSS 0.522594f
C1368 a_n13990_n5465.n108 AVSS 0.792986f
C1369 a_n13990_n5465.t129 AVSS 0.219819f
C1370 a_n13990_n5465.t128 AVSS 0.180853f
C1371 a_n13990_n5465.n109 AVSS 0.636508f
C1372 a_n13990_n5465.n110 AVSS 0.296861f
C1373 a_n13990_n5465.n111 AVSS 2.83331f
C1374 a_n13990_n5465.t137 AVSS 0.522231f
C1375 a_n13990_n5465.t138 AVSS 0.070239f
C1376 a_n13990_n5465.t122 AVSS 0.070239f
C1377 a_n13990_n5465.n112 AVSS 0.275244f
C1378 a_n13990_n5465.n113 AVSS 2.07315f
C1379 a_n13990_n5465.n114 AVSS 9.35673f
C1380 a_n13990_n5465.n115 AVSS 12.59f
C1381 a_n13990_n5465.t80 AVSS 0.073751f
C1382 a_n13990_n5465.t102 AVSS 0.073751f
C1383 a_n13990_n5465.n116 AVSS 0.343286f
C1384 a_n13990_n5465.t48 AVSS 0.333545f
C1385 a_n13990_n5465.t77 AVSS 0.073751f
C1386 a_n13990_n5465.t76 AVSS 0.073751f
C1387 a_n13990_n5465.n117 AVSS 0.343286f
C1388 a_n13990_n5465.t104 AVSS 0.604434f
C1389 a_n13990_n5465.n118 AVSS 1.4001f
C1390 a_n13990_n5465.n119 AVSS 7.42313f
C1391 a_n13990_n5465.n120 AVSS 3.23944f
C1392 a_n13990_n5465.n121 AVSS 0.202914f
C1393 a_n13990_n5465.t97 AVSS 0.073751f
C1394 a_n13990_n5465.t57 AVSS 0.073751f
C1395 a_n13990_n5465.n122 AVSS 0.187146f
C1396 a_n13990_n5465.t96 AVSS 0.073751f
C1397 a_n13990_n5465.t56 AVSS 0.073751f
C1398 a_n13990_n5465.n123 AVSS 0.201973f
C1399 a_n13990_n5465.n124 AVSS 0.512605f
C1400 a_n13990_n5465.n125 AVSS 0.28506f
C1401 a_n13990_n5465.t72 AVSS 0.194302f
C1402 a_n13990_n5465.t71 AVSS 0.20689f
C1403 a_n13990_n5465.n126 AVSS 0.662081f
C1404 a_n13990_n5465.n127 AVSS 0.607929f
C1405 a_n13990_n5465.t47 AVSS 0.194302f
C1406 a_n13990_n5465.t45 AVSS 0.20689f
C1407 a_n13990_n5465.n128 AVSS 0.662081f
C1408 a_n13990_n5465.n129 AVSS 0.607909f
C1409 a_n13990_n5465.t55 AVSS 0.073751f
C1410 a_n13990_n5465.t109 AVSS 0.073751f
C1411 a_n13990_n5465.n130 AVSS 0.187146f
C1412 a_n13990_n5465.t54 AVSS 0.073751f
C1413 a_n13990_n5465.t108 AVSS 0.073751f
C1414 a_n13990_n5465.n131 AVSS 0.201973f
C1415 a_n13990_n5465.n132 AVSS 0.512605f
C1416 a_n13990_n5465.n133 AVSS 0.400355f
C1417 a_n13990_n5465.t33 AVSS 0.194302f
C1418 a_n13990_n5465.t31 AVSS 0.20689f
C1419 a_n13990_n5465.n134 AVSS 0.652343f
C1420 a_n13990_n5465.n135 AVSS 0.597109f
C1421 a_n13990_n5465.t68 AVSS 0.194302f
C1422 a_n13990_n5465.t67 AVSS 0.20689f
C1423 a_n13990_n5465.n136 AVSS 0.655059f
C1424 a_n13990_n5465.n137 AVSS 0.504757f
C1425 a_n13990_n5465.n138 AVSS 0.202914f
C1426 a_n13990_n5465.n139 AVSS 3.23944f
C1427 a_n13990_n5465.t59 AVSS 0.073751f
C1428 a_n13990_n5465.t88 AVSS 0.073751f
C1429 a_n13990_n5465.n140 AVSS 0.708887f
C1430 a_n13990_n5465.t62 AVSS 0.331597f
C1431 a_n13990_n5465.n141 AVSS 1.90188f
C1432 a_n13990_n5465.n142 AVSS 1.40086f
C1433 a_n13990_n5465.t87 AVSS 0.073751f
C1434 a_n13990_n5465.t26 AVSS 0.073751f
C1435 a_n13990_n5465.n143 AVSS 0.340562f
C1436 a_n13990_n5465.n144 AVSS 1.67071f
C1437 a_n13990_n5465.t73 AVSS 0.331597f
C1438 a_n13990_n5465.n145 AVSS 1.09857f
C1439 a_n13990_n5465.n146 AVSS 2.99476f
C1440 a_n13990_n5465.n147 AVSS 3.21714f
C1441 a_n13990_n5465.t28 AVSS 0.073751f
C1442 a_n13990_n5465.t66 AVSS 0.073751f
C1443 a_n13990_n5465.n148 AVSS 0.343286f
C1444 a_n13990_n5465.t30 AVSS 0.333545f
C1445 a_n13990_n5465.t69 AVSS 0.073751f
C1446 a_n13990_n5465.t95 AVSS 0.073751f
C1447 a_n13990_n5465.n149 AVSS 0.343286f
C1448 a_n13990_n5465.t64 AVSS 0.604434f
C1449 a_n13990_n5465.n150 AVSS 1.4001f
C1450 a_n13990_n5465.n151 AVSS 2.79504f
C1451 a_n13990_n5465.n152 AVSS 4.4052f
C1452 a_n13990_n5465.n153 AVSS 0.202914f
C1453 a_n13990_n5465.t58 AVSS 0.194302f
C1454 a_n13990_n5465.t60 AVSS 0.20689f
C1455 a_n13990_n5465.n154 AVSS 0.655059f
C1456 a_n13990_n5465.n155 AVSS 0.504757f
C1457 a_n13990_n5465.n156 AVSS 0.597109f
C1458 a_n13990_n5465.t110 AVSS 0.194302f
C1459 a_n13990_n5465.n157 AVSS 0.652343f
C1460 a_n13990_n5465.t112 AVSS 0.20689f
C1461 VN.t28 AVSS 0.496456f
C1462 VN.n0 AVSS 0.239402f
C1463 VN.n1 AVSS 0.113603f
C1464 VN.n2 AVSS 0.035125f
C1465 VN.n3 AVSS 0.035125f
C1466 VN.n4 AVSS 0.035125f
C1467 VN.n5 AVSS 0.206429f
C1468 VN.n6 AVSS 0.062885f
C1469 VN.t35 AVSS 0.496456f
C1470 VN.n7 AVSS 0.392525f
C1471 VN.n8 AVSS 0.118829f
C1472 VN.n9 AVSS 0.074494f
C1473 VN.n10 AVSS 0.206429f
C1474 VN.n11 AVSS 0.208306f
C1475 VN.t36 AVSS 0.496456f
C1476 VN.n12 AVSS 0.235889f
C1477 VN.n13 AVSS 0.060052f
C1478 VN.n14 AVSS 0.035125f
C1479 VN.n15 AVSS 0.062885f
C1480 VN.n16 AVSS 0.062885f
C1481 VN.n17 AVSS 0.208306f
C1482 VN.n18 AVSS 0.060052f
C1483 VN.t8 AVSS 0.496456f
C1484 VN.n19 AVSS 0.332598f
C1485 VN.n20 AVSS 0.10625f
C1486 VN.n21 AVSS 0.105374f
C1487 VN.n22 AVSS 0.221877f
C1488 VN.n23 AVSS 0.035125f
C1489 VN.n24 AVSS 0.063168f
C1490 VN.n25 AVSS 0.063168f
C1491 VN.n26 AVSS 0.035125f
C1492 VN.n27 AVSS 0.064726f
C1493 VN.n28 AVSS 0.206949f
C1494 VN.n29 AVSS 0.053679f
C1495 VN.t6 AVSS 0.496456f
C1496 VN.n30 AVSS 0.239398f
C1497 VN.n31 AVSS 0.064726f
C1498 VN.n32 AVSS 0.035125f
C1499 VN.n33 AVSS 0.053679f
C1500 VN.n34 AVSS 0.053679f
C1501 VN.n35 AVSS 0.073628f
C1502 VN.t12 AVSS 0.496456f
C1503 VN.n36 AVSS 0.239402f
C1504 VN.n37 AVSS 0.084579f
C1505 VN.n38 AVSS 0.093976f
C1506 VN.n39 AVSS 0.128539f
C1507 VN.n40 AVSS 0.053679f
C1508 VN.n41 AVSS 0.188544f
C1509 VN.n42 AVSS 0.188544f
C1510 VN.n43 AVSS 0.082083f
C1511 VN.n44 AVSS 0.035125f
C1512 VN.n45 AVSS 0.064726f
C1513 VN.n46 AVSS 0.064726f
C1514 VN.n47 AVSS 0.227348f
C1515 VN.n48 AVSS 0.075617f
C1516 VN.t62 AVSS 0.496456f
C1517 VN.n49 AVSS 0.239402f
C1518 VN.n50 AVSS 0.207948f
C1519 VN.n51 AVSS 0.063168f
C1520 VN.n52 AVSS 0.063168f
C1521 VN.n53 AVSS 0.035125f
C1522 VN.n54 AVSS 0.074622f
C1523 VN.t1 AVSS 0.496456f
C1524 VN.n55 AVSS 0.239402f
C1525 VN.n56 AVSS 0.090542f
C1526 VN.n57 AVSS 0.282131f
C1527 VN.n58 AVSS 3.52626f
C1528 VN.n59 AVSS 1.11924f
C1529 VN.n60 AVSS 0.12322f
C1530 VN.n61 AVSS 0.035125f
C1531 VN.n62 AVSS 0.035125f
C1532 VN.n63 AVSS 0.206429f
C1533 VN.n64 AVSS 0.062885f
C1534 VN.t84 AVSS 0.496456f
C1535 VN.n65 AVSS 0.392525f
C1536 VN.n66 AVSS 0.035125f
C1537 VN.n67 AVSS 0.188544f
C1538 VN.n68 AVSS 0.035125f
C1539 VN.n69 AVSS 0.082083f
C1540 VN.n70 AVSS 0.064726f
C1541 VN.n71 AVSS 0.227348f
C1542 VN.t77 AVSS 0.496456f
C1543 VN.n72 AVSS 0.239398f
C1544 VN.n73 AVSS 0.063168f
C1545 VN.t68 AVSS 0.496456f
C1546 VN.n74 AVSS 0.239402f
C1547 VN.n75 AVSS 0.063168f
C1548 VN.n76 AVSS 0.074622f
C1549 VN.n77 AVSS 0.080458f
C1550 VN.t59 AVSS 0.496456f
C1551 VN.n78 AVSS 0.239402f
C1552 VN.n79 AVSS 0.09337f
C1553 VN.n80 AVSS 0.081008f
C1554 VN.n81 AVSS 0.063168f
C1555 VN.n82 AVSS 0.221877f
C1556 VN.n83 AVSS 0.207948f
C1557 VN.n84 AVSS 0.063168f
C1558 VN.n85 AVSS 0.035125f
C1559 VN.n86 AVSS 0.075617f
C1560 VN.n87 AVSS 0.035125f
C1561 VN.n88 AVSS 0.064726f
C1562 VN.n89 AVSS 0.064726f
C1563 VN.n90 AVSS 0.206949f
C1564 VN.n91 AVSS 0.064726f
C1565 VN.n92 AVSS 0.035125f
C1566 VN.n93 AVSS 0.053679f
C1567 VN.n94 AVSS 0.053679f
C1568 VN.n95 AVSS 0.188544f
C1569 VN.n96 AVSS 0.053679f
C1570 VN.n97 AVSS 0.053679f
C1571 VN.n98 AVSS 0.035125f
C1572 VN.n99 AVSS 0.073628f
C1573 VN.t20 AVSS 0.496456f
C1574 VN.n100 AVSS 0.239402f
C1575 VN.n101 AVSS 0.089547f
C1576 VN.n102 AVSS 0.113603f
C1577 VN.n103 AVSS 0.118829f
C1578 VN.n104 AVSS 0.074494f
C1579 VN.n105 AVSS 0.206429f
C1580 VN.n106 AVSS 0.208306f
C1581 VN.t46 AVSS 0.496456f
C1582 VN.n107 AVSS 0.235889f
C1583 VN.n108 AVSS 0.060052f
C1584 VN.n109 AVSS 0.035125f
C1585 VN.n110 AVSS 0.062885f
C1586 VN.n111 AVSS 0.062885f
C1587 VN.n112 AVSS 0.208306f
C1588 VN.n113 AVSS 0.060052f
C1589 VN.t82 AVSS 0.496456f
C1590 VN.n114 AVSS 0.332598f
C1591 VN.n115 AVSS 0.10625f
C1592 VN.n116 AVSS 0.105374f
C1593 VN.n117 AVSS 0.035125f
C1594 VN.n118 AVSS 0.063168f
C1595 VN.n119 AVSS 0.207948f
C1596 VN.n120 AVSS 0.064726f
C1597 VN.t27 AVSS 0.496456f
C1598 VN.n121 AVSS 0.239402f
C1599 VN.n122 AVSS 0.063168f
C1600 VN.n123 AVSS 0.035125f
C1601 VN.n124 AVSS 0.064726f
C1602 VN.n125 AVSS 0.064726f
C1603 VN.t73 AVSS 0.496456f
C1604 VN.n126 AVSS 0.239398f
C1605 VN.n127 AVSS 0.053679f
C1606 VN.n128 AVSS 0.035125f
C1607 VN.n129 AVSS 0.053679f
C1608 VN.n130 AVSS 0.053679f
C1609 VN.n131 AVSS 0.073628f
C1610 VN.n132 AVSS 0.39827f
C1611 VN.t63 AVSS 0.496456f
C1612 VN.n133 AVSS 0.239402f
C1613 VN.n134 AVSS 0.035125f
C1614 VN.n135 AVSS 0.035125f
C1615 VN.n136 AVSS 0.221877f
C1616 VN.n137 AVSS 0.035125f
C1617 VN.n138 AVSS 0.063168f
C1618 VN.n139 AVSS 0.063168f
C1619 VN.n140 AVSS 0.035125f
C1620 VN.n141 AVSS 0.064726f
C1621 VN.n142 AVSS 0.206949f
C1622 VN.n143 AVSS 0.053679f
C1623 VN.t30 AVSS 0.496456f
C1624 VN.n144 AVSS 0.239398f
C1625 VN.n145 AVSS 0.064726f
C1626 VN.n146 AVSS 0.035125f
C1627 VN.n147 AVSS 0.053679f
C1628 VN.n148 AVSS 0.053679f
C1629 VN.n149 AVSS 0.073628f
C1630 VN.n150 AVSS 0.120455f
C1631 VN.n151 AVSS 0.035125f
C1632 VN.n152 AVSS 0.048753f
C1633 VN.n153 AVSS 0.035125f
C1634 VN.n154 AVSS 0.218893f
C1635 VN.n155 AVSS 0.062885f
C1636 VN.t19 AVSS 0.496456f
C1637 VN.n156 AVSS 0.405555f
C1638 VN.n157 AVSS 0.035125f
C1639 VN.n158 AVSS 0.061688f
C1640 VN.n159 AVSS 0.062885f
C1641 VN.n160 AVSS 0.149241f
C1642 VN.n161 AVSS 0.064726f
C1643 VN.n162 AVSS 0.061684f
C1644 VN.n163 AVSS 0.062885f
C1645 VN.n164 AVSS 0.061688f
C1646 VN.n165 AVSS 0.063168f
C1647 VN.n166 AVSS 0.061688f
C1648 VN.n167 AVSS 0.062885f
C1649 VN.n168 AVSS 0.061688f
C1650 VN.n169 AVSS 0.39827f
C1651 VN.n170 AVSS 0.116294f
C1652 VN.n171 AVSS 0.035125f
C1653 VN.t66 AVSS 0.496456f
C1654 VN.n172 AVSS 0.229452f
C1655 VN.n173 AVSS 0.053679f
C1656 VN.n174 AVSS 0.136806f
C1657 VN.n175 AVSS 0.035125f
C1658 VN.n176 AVSS 0.059694f
C1659 VN.n177 AVSS 0.064726f
C1660 VN.n178 AVSS 0.159195f
C1661 VN.n179 AVSS 0.035125f
C1662 VN.t29 AVSS 0.496456f
C1663 VN.n180 AVSS 0.193633f
C1664 VN.n181 AVSS 0.063168f
C1665 VN.n182 AVSS 0.159195f
C1666 VN.n183 AVSS 0.035125f
C1667 VN.t34 AVSS 0.496456f
C1668 VN.n184 AVSS 0.192638f
C1669 VN.n185 AVSS 0.035125f
C1670 VN.n186 AVSS 0.218893f
C1671 VN.n187 AVSS 0.062885f
C1672 VN.t51 AVSS 0.496456f
C1673 VN.n188 AVSS 0.405555f
C1674 VN.n189 AVSS 0.035125f
C1675 VN.t21 AVSS 0.496456f
C1676 VN.n190 AVSS 0.229452f
C1677 VN.n191 AVSS 0.062885f
C1678 VN.n192 AVSS 0.149241f
C1679 VN.n193 AVSS 0.064726f
C1680 VN.t78 AVSS 0.496456f
C1681 VN.n194 AVSS 0.200099f
C1682 VN.n195 AVSS 0.062885f
C1683 VN.n196 AVSS 0.061688f
C1684 VN.n197 AVSS 0.063168f
C1685 VN.n198 AVSS 0.061688f
C1686 VN.n199 AVSS 0.131563f
C1687 VN.n200 AVSS 0.061688f
C1688 VN.n201 AVSS 0.126444f
C1689 VN.t60 AVSS 0.496456f
C1690 VN.n202 AVSS 0.237615f
C1691 VN.n203 AVSS 0.059698f
C1692 VN.n204 AVSS 0.08086f
C1693 VN.n205 AVSS 0.063168f
C1694 VN.n206 AVSS 0.159195f
C1695 VN.n207 AVSS 0.16019f
C1696 VN.n208 AVSS 0.062885f
C1697 VN.n209 AVSS 0.062885f
C1698 VN.n210 AVSS 0.035125f
C1699 VN.n211 AVSS 0.047758f
C1700 VN.t70 AVSS 0.496456f
C1701 VN.n212 AVSS 0.193633f
C1702 VN.n213 AVSS 0.059698f
C1703 VN.n214 AVSS 0.035125f
C1704 VN.n215 AVSS 0.064726f
C1705 VN.n216 AVSS 0.159195f
C1706 VN.n217 AVSS 0.16566f
C1707 VN.n218 AVSS 0.061684f
C1708 VN.n219 AVSS 0.041289f
C1709 VN.n220 AVSS 0.035125f
C1710 VN.n221 AVSS 0.062885f
C1711 VN.n222 AVSS 0.061684f
C1712 VN.n223 AVSS 0.059694f
C1713 VN.n224 AVSS 0.035125f
C1714 VN.n225 AVSS 0.053679f
C1715 VN.n226 AVSS 0.053679f
C1716 VN.n227 AVSS 0.136806f
C1717 VN.n228 AVSS 0.061688f
C1718 VN.n229 AVSS 0.061688f
C1719 VN.n230 AVSS 0.01194f
C1720 VN.n231 AVSS 0.035125f
C1721 VN.n232 AVSS 0.120455f
C1722 VN.n233 AVSS 0.107388f
C1723 VN.n234 AVSS 0.1136f
C1724 VN.n235 AVSS 0.11883f
C1725 VN.n236 AVSS 0.074496f
C1726 VN.n237 AVSS 0.218893f
C1727 VN.n238 AVSS 0.220882f
C1728 VN.t42 AVSS 0.496456f
C1729 VN.n239 AVSS 0.239402f
C1730 VN.n240 AVSS 0.063678f
C1731 VN.n241 AVSS 0.035125f
C1732 VN.n242 AVSS 0.062885f
C1733 VN.n243 AVSS 0.062885f
C1734 VN.n244 AVSS 0.220882f
C1735 VN.n245 AVSS 0.063678f
C1736 VN.t69 AVSS 0.496456f
C1737 VN.n246 AVSS 0.342002f
C1738 VN.n247 AVSS 0.106251f
C1739 VN.n248 AVSS 0.277999f
C1740 VN.n249 AVSS 0.048753f
C1741 VN.n250 AVSS 0.116294f
C1742 VN.n251 AVSS 0.105374f
C1743 VN.n252 AVSS 0.035125f
C1744 VN.n253 AVSS 0.059698f
C1745 VN.n254 AVSS 0.061688f
C1746 VN.n255 AVSS 0.062885f
C1747 VN.n256 AVSS 0.062885f
C1748 VN.n257 AVSS 0.16019f
C1749 VN.n258 AVSS 0.047758f
C1750 VN.n259 AVSS 0.061688f
C1751 VN.n260 AVSS 0.063168f
C1752 VN.n261 AVSS 0.035125f
C1753 VN.n262 AVSS 0.059698f
C1754 VN.n263 AVSS 0.061688f
C1755 VN.n264 AVSS 0.062885f
C1756 VN.n265 AVSS 0.062885f
C1757 VN.n266 AVSS 0.16566f
C1758 VN.t75 AVSS 0.496456f
C1759 VN.n267 AVSS 0.200099f
C1760 VN.n268 AVSS 0.041289f
C1761 VN.n269 AVSS 0.061684f
C1762 VN.n270 AVSS 0.064726f
C1763 VN.n271 AVSS 0.035125f
C1764 VN.n272 AVSS 0.053679f
C1765 VN.n273 AVSS 0.149241f
C1766 VN.n274 AVSS 0.061684f
C1767 VN.n275 AVSS 0.062885f
C1768 VN.n276 AVSS 0.062885f
C1769 VN.n277 AVSS 0.061688f
C1770 VN.n278 AVSS 0.01194f
C1771 VN.n279 AVSS 0.061688f
C1772 VN.n280 AVSS 0.035125f
C1773 VN.n281 AVSS 0.39827f
C1774 VN.n282 AVSS 0.112356f
C1775 VN.n283 AVSS 0.391263f
C1776 VN.n284 AVSS 0.391305f
C1777 VN.n285 AVSS 0.035125f
C1778 VN.n286 AVSS 0.048753f
C1779 VN.t72 AVSS 0.496456f
C1780 VN.n287 AVSS 0.192638f
C1781 VN.n288 AVSS 0.059698f
C1782 VN.n289 AVSS 0.035125f
C1783 VN.n290 AVSS 0.063168f
C1784 VN.n291 AVSS 0.159195f
C1785 VN.n292 AVSS 0.16019f
C1786 VN.n293 AVSS 0.062885f
C1787 VN.n294 AVSS 0.035125f
C1788 VN.n295 AVSS 0.047758f
C1789 VN.t11 AVSS 0.496456f
C1790 VN.n296 AVSS 0.193633f
C1791 VN.n297 AVSS 0.059698f
C1792 VN.n298 AVSS 0.035125f
C1793 VN.n299 AVSS 0.064726f
C1794 VN.n300 AVSS 0.159195f
C1795 VN.n301 AVSS 0.16566f
C1796 VN.n302 AVSS 0.062885f
C1797 VN.n303 AVSS 0.035125f
C1798 VN.n304 AVSS 0.041289f
C1799 VN.t31 AVSS 0.496456f
C1800 VN.n305 AVSS 0.200099f
C1801 VN.n306 AVSS 0.061684f
C1802 VN.n307 AVSS 0.059694f
C1803 VN.n308 AVSS 0.035125f
C1804 VN.n309 AVSS 0.053679f
C1805 VN.n310 AVSS 0.053679f
C1806 VN.n311 AVSS 0.136806f
C1807 VN.n312 AVSS 0.061688f
C1808 VN.n313 AVSS 0.062885f
C1809 VN.n314 AVSS 0.035125f
C1810 VN.n315 AVSS 0.01194f
C1811 VN.t54 AVSS 0.496456f
C1812 VN.n316 AVSS 0.229452f
C1813 VN.n317 AVSS 0.107388f
C1814 VN.n318 AVSS 0.1136f
C1815 VN.n319 AVSS 0.11883f
C1816 VN.n320 AVSS 0.074496f
C1817 VN.n321 AVSS 0.218893f
C1818 VN.n322 AVSS 0.220882f
C1819 VN.t80 AVSS 0.496456f
C1820 VN.n323 AVSS 0.239402f
C1821 VN.n324 AVSS 0.063678f
C1822 VN.n325 AVSS 0.035125f
C1823 VN.n326 AVSS 0.062885f
C1824 VN.n327 AVSS 0.062885f
C1825 VN.n328 AVSS 0.220882f
C1826 VN.n329 AVSS 0.063678f
C1827 VN.t18 AVSS 0.496456f
C1828 VN.n330 AVSS 0.342002f
C1829 VN.n331 AVSS 0.106251f
C1830 VN.n332 AVSS 0.063168f
C1831 VN.t2 AVSS 0.496456f
C1832 VN.n333 AVSS 0.192638f
C1833 VN.n334 AVSS 0.159195f
C1834 VN.n335 AVSS 0.035125f
C1835 VN.n336 AVSS 0.047758f
C1836 VN.n337 AVSS 0.064726f
C1837 VN.t85 AVSS 0.496456f
C1838 VN.n338 AVSS 0.193633f
C1839 VN.n339 AVSS 0.159195f
C1840 VN.n340 AVSS 0.035125f
C1841 VN.n341 AVSS 0.041289f
C1842 VN.n342 AVSS 0.053679f
C1843 VN.t38 AVSS 0.496456f
C1844 VN.n343 AVSS 0.200099f
C1845 VN.n344 AVSS 0.149241f
C1846 VN.n345 AVSS 0.079159f
C1847 VN.n346 AVSS 0.136806f
C1848 VN.n347 AVSS 0.01194f
C1849 VN.n348 AVSS 0.053679f
C1850 VN.t14 AVSS 0.496456f
C1851 VN.n349 AVSS 0.229452f
C1852 VN.n350 AVSS 0.116615f
C1853 VN.n351 AVSS 0.128539f
C1854 VN.n352 AVSS 0.061688f
C1855 VN.n353 AVSS 0.061688f
C1856 VN.n354 AVSS 0.062885f
C1857 VN.n355 AVSS 0.062885f
C1858 VN.n356 AVSS 0.061684f
C1859 VN.n357 AVSS 0.059694f
C1860 VN.n358 AVSS 0.035125f
C1861 VN.n359 AVSS 0.064726f
C1862 VN.n360 AVSS 0.061684f
C1863 VN.n361 AVSS 0.16566f
C1864 VN.n362 AVSS 0.062885f
C1865 VN.n363 AVSS 0.062885f
C1866 VN.n364 AVSS 0.061688f
C1867 VN.n365 AVSS 0.059698f
C1868 VN.n366 AVSS 0.035125f
C1869 VN.n367 AVSS 0.063168f
C1870 VN.n368 AVSS 0.061688f
C1871 VN.n369 AVSS 0.16019f
C1872 VN.n370 AVSS 0.062885f
C1873 VN.n371 AVSS 0.062885f
C1874 VN.n372 AVSS 0.061688f
C1875 VN.n373 AVSS 0.059698f
C1876 VN.n374 AVSS 0.035125f
C1877 VN.n375 AVSS 0.105374f
C1878 VN.n376 AVSS 0.116294f
C1879 VN.n377 AVSS 0.277999f
C1880 VN.n378 AVSS 1.11924f
C1881 VN.n379 AVSS 5.51141f
C1882 VN.n380 AVSS 0.370227f
C1883 VN.t52 AVSS 0.496456f
C1884 VN.n381 AVSS 0.239402f
C1885 VN.n382 AVSS 0.035125f
C1886 VN.n383 AVSS 0.074494f
C1887 VN.n384 AVSS 0.060052f
C1888 VN.n385 AVSS 0.062885f
C1889 VN.t17 AVSS 0.496456f
C1890 VN.n386 AVSS 0.235889f
C1891 VN.t48 AVSS 0.496456f
C1892 VN.n387 AVSS 0.332598f
C1893 VN.n388 AVSS 0.035125f
C1894 VN.t0 AVSS 0.496456f
C1895 VN.n389 AVSS 0.239402f
C1896 VN.n390 AVSS 0.063168f
C1897 VN.n391 AVSS 0.063168f
C1898 VN.n392 AVSS 0.063168f
C1899 VN.t83 AVSS 0.496456f
C1900 VN.n393 AVSS 0.239402f
C1901 VN.n394 AVSS 0.064726f
C1902 VN.n395 AVSS 0.035125f
C1903 VN.n396 AVSS 0.064726f
C1904 VN.n397 AVSS 0.064726f
C1905 VN.t37 AVSS 0.496456f
C1906 VN.n398 AVSS 0.239398f
C1907 VN.n399 AVSS 0.053679f
C1908 VN.n400 AVSS 0.035125f
C1909 VN.n401 AVSS 0.053679f
C1910 VN.n402 AVSS 0.053679f
C1911 VN.n403 AVSS 0.073628f
C1912 VN.t13 AVSS 0.496456f
C1913 VN.n404 AVSS 0.239402f
C1914 VN.n405 AVSS 0.128539f
C1915 VN.n406 AVSS 0.093976f
C1916 VN.n407 AVSS 0.084579f
C1917 VN.n408 AVSS 0.053679f
C1918 VN.n409 AVSS 0.188544f
C1919 VN.n410 AVSS 0.188544f
C1920 VN.n411 AVSS 0.082083f
C1921 VN.n412 AVSS 0.035125f
C1922 VN.n413 AVSS 0.064726f
C1923 VN.n414 AVSS 0.206949f
C1924 VN.n415 AVSS 0.227348f
C1925 VN.n416 AVSS 0.075617f
C1926 VN.n417 AVSS 0.035125f
C1927 VN.n418 AVSS 0.063168f
C1928 VN.n419 AVSS 0.207948f
C1929 VN.n420 AVSS 0.221877f
C1930 VN.n421 AVSS 0.074622f
C1931 VN.n422 AVSS 0.035125f
C1932 VN.n423 AVSS 0.282131f
C1933 VN.n424 AVSS 0.090542f
C1934 VN.n425 AVSS 0.105374f
C1935 VN.n426 AVSS 0.10625f
C1936 VN.n427 AVSS 0.035125f
C1937 VN.n428 AVSS 0.060052f
C1938 VN.n429 AVSS 0.208306f
C1939 VN.n430 AVSS 0.206429f
C1940 VN.n431 AVSS 0.062885f
C1941 VN.n432 AVSS 0.035125f
C1942 VN.n433 AVSS 0.062885f
C1943 VN.n434 AVSS 0.208306f
C1944 VN.n435 AVSS 0.206429f
C1945 VN.t43 AVSS 0.496456f
C1946 VN.n436 AVSS 0.392525f
C1947 VN.n437 AVSS 0.118829f
C1948 VN.n438 AVSS 0.113603f
C1949 VN.n439 AVSS 0.089547f
C1950 VN.n440 AVSS 0.12322f
C1951 VN.n441 AVSS 0.035125f
C1952 VN.n442 AVSS 0.053679f
C1953 VN.n443 AVSS 0.188544f
C1954 VN.n444 AVSS 0.188544f
C1955 VN.n445 AVSS 0.082083f
C1956 VN.n446 AVSS 0.035125f
C1957 VN.n447 AVSS 0.064726f
C1958 VN.n448 AVSS 0.064726f
C1959 VN.n449 AVSS 0.227348f
C1960 VN.n450 AVSS 0.075617f
C1961 VN.t7 AVSS 0.496456f
C1962 VN.n451 AVSS 0.239402f
C1963 VN.n452 AVSS 0.207948f
C1964 VN.n453 AVSS 0.063168f
C1965 VN.n454 AVSS 0.063168f
C1966 VN.n455 AVSS 0.035125f
C1967 VN.n456 AVSS 0.074622f
C1968 VN.t71 AVSS 0.496456f
C1969 VN.n457 AVSS 0.239402f
C1970 VN.n458 AVSS 0.090542f
C1971 VN.n459 AVSS 0.39827f
C1972 VN.n460 AVSS 0.39827f
C1973 VN.n461 AVSS 0.089547f
C1974 VN.n462 AVSS 0.39827f
C1975 VN.n463 AVSS 0.035125f
C1976 VN.n464 AVSS 0.053679f
C1977 VN.n465 AVSS 0.188544f
C1978 VN.n466 AVSS 0.188544f
C1979 VN.n467 AVSS 0.082083f
C1980 VN.n468 AVSS 0.035125f
C1981 VN.n469 AVSS 0.064726f
C1982 VN.n470 AVSS 0.206949f
C1983 VN.n471 AVSS 0.227348f
C1984 VN.n472 AVSS 0.075617f
C1985 VN.n473 AVSS 0.035125f
C1986 VN.n474 AVSS 0.063168f
C1987 VN.n475 AVSS 0.063168f
C1988 VN.n476 AVSS 0.221877f
C1989 VN.n477 AVSS 0.074622f
C1990 VN.t33 AVSS 0.496456f
C1991 VN.n478 AVSS 0.239402f
C1992 VN.n479 AVSS 0.090542f
C1993 VN.n480 AVSS 0.282131f
C1994 VN.n481 AVSS 0.370227f
C1995 VN.n482 AVSS 5.51141f
C1996 VN.n483 AVSS 0.120455f
C1997 VN.n484 AVSS 0.035125f
C1998 VN.n485 AVSS 0.048753f
C1999 VN.n486 AVSS 0.035125f
C2000 VN.n487 AVSS 0.218893f
C2001 VN.n488 AVSS 0.062885f
C2002 VN.t39 AVSS 0.496456f
C2003 VN.n489 AVSS 0.405555f
C2004 VN.n490 AVSS 0.035125f
C2005 VN.n491 AVSS 0.061688f
C2006 VN.n492 AVSS 0.062885f
C2007 VN.n493 AVSS 0.149241f
C2008 VN.n494 AVSS 0.064726f
C2009 VN.n495 AVSS 0.061684f
C2010 VN.n496 AVSS 0.062885f
C2011 VN.n497 AVSS 0.061688f
C2012 VN.n498 AVSS 0.063168f
C2013 VN.n499 AVSS 0.061688f
C2014 VN.n500 AVSS 0.131563f
C2015 VN.n501 AVSS 0.061688f
C2016 VN.n502 AVSS 0.126444f
C2017 VN.t74 AVSS 0.496456f
C2018 VN.n503 AVSS 0.237615f
C2019 VN.n504 AVSS 0.059698f
C2020 VN.n505 AVSS 0.08086f
C2021 VN.n506 AVSS 0.063168f
C2022 VN.n507 AVSS 0.159195f
C2023 VN.n508 AVSS 0.16019f
C2024 VN.n509 AVSS 0.062885f
C2025 VN.n510 AVSS 0.035125f
C2026 VN.n511 AVSS 0.047758f
C2027 VN.t22 AVSS 0.496456f
C2028 VN.n512 AVSS 0.193633f
C2029 VN.n513 AVSS 0.059698f
C2030 VN.n514 AVSS 0.035125f
C2031 VN.n515 AVSS 0.064726f
C2032 VN.n516 AVSS 0.159195f
C2033 VN.n517 AVSS 0.16566f
C2034 VN.n518 AVSS 0.062885f
C2035 VN.n519 AVSS 0.035125f
C2036 VN.n520 AVSS 0.041289f
C2037 VN.t47 AVSS 0.496456f
C2038 VN.n521 AVSS 0.200099f
C2039 VN.n522 AVSS 0.061684f
C2040 VN.n523 AVSS 0.059694f
C2041 VN.n524 AVSS 0.035125f
C2042 VN.n525 AVSS 0.053679f
C2043 VN.n526 AVSS 0.053679f
C2044 VN.n527 AVSS 0.136806f
C2045 VN.n528 AVSS 0.061688f
C2046 VN.n529 AVSS 0.062885f
C2047 VN.n530 AVSS 0.035125f
C2048 VN.n531 AVSS 0.01194f
C2049 VN.t44 AVSS 0.496456f
C2050 VN.n532 AVSS 0.229452f
C2051 VN.n533 AVSS 0.107388f
C2052 VN.n534 AVSS 0.1136f
C2053 VN.n535 AVSS 0.11883f
C2054 VN.n536 AVSS 0.074496f
C2055 VN.n537 AVSS 0.218893f
C2056 VN.n538 AVSS 0.220882f
C2057 VN.t25 AVSS 0.496456f
C2058 VN.n539 AVSS 0.239402f
C2059 VN.n540 AVSS 0.063678f
C2060 VN.n541 AVSS 0.035125f
C2061 VN.n542 AVSS 0.062885f
C2062 VN.n543 AVSS 0.062885f
C2063 VN.n544 AVSS 0.220882f
C2064 VN.n545 AVSS 0.063678f
C2065 VN.t86 AVSS 0.496456f
C2066 VN.n546 AVSS 0.342002f
C2067 VN.n547 AVSS 0.106251f
C2068 VN.n548 AVSS 0.063168f
C2069 VN.t79 AVSS 0.496456f
C2070 VN.n549 AVSS 0.192638f
C2071 VN.n550 AVSS 0.159195f
C2072 VN.n551 AVSS 0.035125f
C2073 VN.n552 AVSS 0.047758f
C2074 VN.n553 AVSS 0.064726f
C2075 VN.t57 AVSS 0.496456f
C2076 VN.n554 AVSS 0.193633f
C2077 VN.n555 AVSS 0.159195f
C2078 VN.n556 AVSS 0.035125f
C2079 VN.n557 AVSS 0.041289f
C2080 VN.n558 AVSS 0.053679f
C2081 VN.t3 AVSS 0.496456f
C2082 VN.n559 AVSS 0.200099f
C2083 VN.n560 AVSS 0.149241f
C2084 VN.n561 AVSS 0.035125f
C2085 VN.n562 AVSS 0.136806f
C2086 VN.n563 AVSS 0.01194f
C2087 VN.n564 AVSS 0.053679f
C2088 VN.n565 AVSS 0.39827f
C2089 VN.t65 AVSS 0.496456f
C2090 VN.n566 AVSS 0.229452f
C2091 VN.n567 AVSS 0.035125f
C2092 VN.n568 AVSS 0.061688f
C2093 VN.n569 AVSS 0.063168f
C2094 VN.n570 AVSS 0.061688f
C2095 VN.n571 AVSS 0.062885f
C2096 VN.n572 AVSS 0.062885f
C2097 VN.n573 AVSS 0.061688f
C2098 VN.n574 AVSS 0.064726f
C2099 VN.n575 AVSS 0.061684f
C2100 VN.n576 AVSS 0.062885f
C2101 VN.n577 AVSS 0.061684f
C2102 VN.n578 AVSS 0.053679f
C2103 VN.n579 AVSS 0.061688f
C2104 VN.n580 AVSS 0.120455f
C2105 VN.n581 AVSS 0.035125f
C2106 VN.n582 AVSS 0.074496f
C2107 VN.n583 AVSS 0.063678f
C2108 VN.n584 AVSS 0.062885f
C2109 VN.t53 AVSS 0.496456f
C2110 VN.n585 AVSS 0.239402f
C2111 VN.t24 AVSS 0.496456f
C2112 VN.n586 AVSS 0.342002f
C2113 VN.n587 AVSS 0.035125f
C2114 VN.n588 AVSS 0.363145f
C2115 VN.n589 AVSS 0.277999f
C2116 VN.t87 AVSS 0.496456f
C2117 VN.n590 AVSS 0.192638f
C2118 VN.n591 AVSS 0.062885f
C2119 VN.n592 AVSS 0.059698f
C2120 VN.n593 AVSS 0.16019f
C2121 VN.n594 AVSS 0.035125f
C2122 VN.t61 AVSS 0.496456f
C2123 VN.n595 AVSS 0.193633f
C2124 VN.n596 AVSS 0.062885f
C2125 VN.n597 AVSS 0.059698f
C2126 VN.n598 AVSS 0.16566f
C2127 VN.n599 AVSS 0.035125f
C2128 VN.t5 AVSS 0.496456f
C2129 VN.n600 AVSS 0.200099f
C2130 VN.n601 AVSS 0.062885f
C2131 VN.n602 AVSS 0.059694f
C2132 VN.n603 AVSS 0.136806f
C2133 VN.n604 AVSS 0.116615f
C2134 VN.n605 AVSS 0.061688f
C2135 VN.t9 AVSS 0.496456f
C2136 VN.n606 AVSS 0.229452f
C2137 VN.n607 AVSS 0.079159f
C2138 VN.n608 AVSS 0.01194f
C2139 VN.n609 AVSS 0.061688f
C2140 VN.n610 AVSS 0.128539f
C2141 VN.n611 AVSS 0.053679f
C2142 VN.n612 AVSS 0.053679f
C2143 VN.n613 AVSS 0.149241f
C2144 VN.n614 AVSS 0.061684f
C2145 VN.n615 AVSS 0.062885f
C2146 VN.n616 AVSS 0.035125f
C2147 VN.n617 AVSS 0.041289f
C2148 VN.n618 AVSS 0.061684f
C2149 VN.n619 AVSS 0.064726f
C2150 VN.n620 AVSS 0.064726f
C2151 VN.n621 AVSS 0.159195f
C2152 VN.n622 AVSS 0.061688f
C2153 VN.n623 AVSS 0.062885f
C2154 VN.n624 AVSS 0.035125f
C2155 VN.n625 AVSS 0.047758f
C2156 VN.n626 AVSS 0.061688f
C2157 VN.n627 AVSS 0.063168f
C2158 VN.n628 AVSS 0.063168f
C2159 VN.n629 AVSS 0.159195f
C2160 VN.n630 AVSS 0.061688f
C2161 VN.n631 AVSS 0.062885f
C2162 VN.n632 AVSS 0.035125f
C2163 VN.n633 AVSS 0.048753f
C2164 VN.n634 AVSS 0.116294f
C2165 VN.n635 AVSS 0.105374f
C2166 VN.n636 AVSS 0.106251f
C2167 VN.n637 AVSS 0.035125f
C2168 VN.n638 AVSS 0.063678f
C2169 VN.n639 AVSS 0.220882f
C2170 VN.n640 AVSS 0.218893f
C2171 VN.n641 AVSS 0.062885f
C2172 VN.n642 AVSS 0.035125f
C2173 VN.n643 AVSS 0.062885f
C2174 VN.n644 AVSS 0.220882f
C2175 VN.n645 AVSS 0.218893f
C2176 VN.t50 AVSS 0.496456f
C2177 VN.n646 AVSS 0.405555f
C2178 VN.n647 AVSS 0.11883f
C2179 VN.n648 AVSS 0.1136f
C2180 VN.n649 AVSS 0.107388f
C2181 VN.t26 AVSS 0.496456f
C2182 VN.n650 AVSS 0.229452f
C2183 VN.n651 AVSS 0.01194f
C2184 VN.n652 AVSS 0.035125f
C2185 VN.n653 AVSS 0.062885f
C2186 VN.n654 AVSS 0.061688f
C2187 VN.n655 AVSS 0.136806f
C2188 VN.n656 AVSS 0.149241f
C2189 VN.n657 AVSS 0.053679f
C2190 VN.n658 AVSS 0.035125f
C2191 VN.n659 AVSS 0.059694f
C2192 VN.t55 AVSS 0.496456f
C2193 VN.n660 AVSS 0.200099f
C2194 VN.n661 AVSS 0.041289f
C2195 VN.n662 AVSS 0.035125f
C2196 VN.n663 AVSS 0.062885f
C2197 VN.n664 AVSS 0.16566f
C2198 VN.n665 AVSS 0.159195f
C2199 VN.n666 AVSS 0.064726f
C2200 VN.n667 AVSS 0.035125f
C2201 VN.n668 AVSS 0.059698f
C2202 VN.t15 AVSS 0.496456f
C2203 VN.n669 AVSS 0.193633f
C2204 VN.n670 AVSS 0.047758f
C2205 VN.n671 AVSS 0.035125f
C2206 VN.n672 AVSS 0.062885f
C2207 VN.n673 AVSS 0.16019f
C2208 VN.n674 AVSS 0.159195f
C2209 VN.n675 AVSS 0.063168f
C2210 VN.n676 AVSS 0.035125f
C2211 VN.n677 AVSS 0.059698f
C2212 VN.t40 AVSS 0.496456f
C2213 VN.n678 AVSS 0.192638f
C2214 VN.n679 AVSS 0.048753f
C2215 VN.n680 AVSS 0.116294f
C2216 VN.n681 AVSS 0.391305f
C2217 VN.n682 AVSS 0.391263f
C2218 VN.n683 AVSS 0.112356f
C2219 VN.n684 AVSS 0.39827f
C2220 VN.n685 AVSS 0.035125f
C2221 VN.n686 AVSS 0.061688f
C2222 VN.n687 AVSS 0.061688f
C2223 VN.n688 AVSS 0.062885f
C2224 VN.n689 AVSS 0.062885f
C2225 VN.n690 AVSS 0.061684f
C2226 VN.n691 AVSS 0.059694f
C2227 VN.n692 AVSS 0.035125f
C2228 VN.n693 AVSS 0.064726f
C2229 VN.n694 AVSS 0.061684f
C2230 VN.n695 AVSS 0.16566f
C2231 VN.n696 AVSS 0.062885f
C2232 VN.n697 AVSS 0.062885f
C2233 VN.n698 AVSS 0.061688f
C2234 VN.n699 AVSS 0.059698f
C2235 VN.n700 AVSS 0.035125f
C2236 VN.n701 AVSS 0.063168f
C2237 VN.n702 AVSS 0.061688f
C2238 VN.n703 AVSS 0.16019f
C2239 VN.n704 AVSS 0.062885f
C2240 VN.n705 AVSS 0.062885f
C2241 VN.n706 AVSS 0.061688f
C2242 VN.n707 AVSS 0.059698f
C2243 VN.n708 AVSS 0.035125f
C2244 VN.n709 AVSS 0.105374f
C2245 VN.n710 AVSS 0.116294f
C2246 VN.n711 AVSS 0.277999f
C2247 VN.n712 AVSS 0.363145f
C2248 VN.n713 AVSS 3.52626f
C2249 VN.n714 AVSS 0.12322f
C2250 VN.n715 AVSS 0.035125f
C2251 VN.n716 AVSS 0.035125f
C2252 VN.n717 AVSS 0.206429f
C2253 VN.n718 AVSS 0.062885f
C2254 VN.t32 AVSS 0.496456f
C2255 VN.n719 AVSS 0.392525f
C2256 VN.n720 AVSS 0.035125f
C2257 VN.n721 AVSS 0.188544f
C2258 VN.n722 AVSS 0.035125f
C2259 VN.n723 AVSS 0.082083f
C2260 VN.n724 AVSS 0.064726f
C2261 VN.n725 AVSS 0.227348f
C2262 VN.n726 AVSS 0.063168f
C2263 VN.t23 AVSS 0.496456f
C2264 VN.n727 AVSS 0.239402f
C2265 VN.n728 AVSS 0.063168f
C2266 VN.n729 AVSS 0.074622f
C2267 VN.t76 AVSS 0.496456f
C2268 VN.n730 AVSS 0.239402f
C2269 VN.n731 AVSS 0.080458f
C2270 VN.n732 AVSS 0.09337f
C2271 VN.n733 AVSS 0.081008f
C2272 VN.n734 AVSS 0.063168f
C2273 VN.n735 AVSS 0.221877f
C2274 VN.n736 AVSS 0.207948f
C2275 VN.n737 AVSS 0.063168f
C2276 VN.n738 AVSS 0.035125f
C2277 VN.n739 AVSS 0.075617f
C2278 VN.n740 AVSS 0.035125f
C2279 VN.n741 AVSS 0.064726f
C2280 VN.n742 AVSS 0.064726f
C2281 VN.t49 AVSS 0.496456f
C2282 VN.n743 AVSS 0.239398f
C2283 VN.n744 AVSS 0.206949f
C2284 VN.n745 AVSS 0.064726f
C2285 VN.n746 AVSS 0.035125f
C2286 VN.n747 AVSS 0.053679f
C2287 VN.n748 AVSS 0.053679f
C2288 VN.n749 AVSS 0.188544f
C2289 VN.n750 AVSS 0.053679f
C2290 VN.n751 AVSS 0.053679f
C2291 VN.n752 AVSS 0.035125f
C2292 VN.n753 AVSS 0.073628f
C2293 VN.t45 AVSS 0.496456f
C2294 VN.n754 AVSS 0.239402f
C2295 VN.n755 AVSS 0.089547f
C2296 VN.n756 AVSS 0.113603f
C2297 VN.n757 AVSS 0.118829f
C2298 VN.n758 AVSS 0.074494f
C2299 VN.n759 AVSS 0.206429f
C2300 VN.n760 AVSS 0.208306f
C2301 VN.t10 AVSS 0.496456f
C2302 VN.n761 AVSS 0.235889f
C2303 VN.n762 AVSS 0.060052f
C2304 VN.n763 AVSS 0.035125f
C2305 VN.n764 AVSS 0.062885f
C2306 VN.n765 AVSS 0.062885f
C2307 VN.n766 AVSS 0.208306f
C2308 VN.n767 AVSS 0.060052f
C2309 VN.t64 AVSS 0.496456f
C2310 VN.n768 AVSS 0.332598f
C2311 VN.n769 AVSS 0.10625f
C2312 VN.n770 AVSS 0.105374f
C2313 VN.n771 AVSS 0.221877f
C2314 VN.n772 AVSS 0.035125f
C2315 VN.n773 AVSS 0.063168f
C2316 VN.n774 AVSS 0.063168f
C2317 VN.n775 AVSS 0.035125f
C2318 VN.n776 AVSS 0.064726f
C2319 VN.n777 AVSS 0.206949f
C2320 VN.n778 AVSS 0.053679f
C2321 VN.t4 AVSS 0.496456f
C2322 VN.n779 AVSS 0.239398f
C2323 VN.n780 AVSS 0.064726f
C2324 VN.n781 AVSS 0.035125f
C2325 VN.n782 AVSS 0.053679f
C2326 VN.n783 AVSS 0.053679f
C2327 VN.n784 AVSS 0.073628f
C2328 VN.n785 AVSS 0.39827f
C2329 VN.t67 AVSS 0.496456f
C2330 VN.n786 AVSS 0.239402f
C2331 VN.n787 AVSS 0.035125f
C2332 VN.n788 AVSS 0.035125f
C2333 VN.n789 AVSS 0.035125f
C2334 VN.n790 AVSS 0.063168f
C2335 VN.n791 AVSS 0.207948f
C2336 VN.n792 AVSS 0.064726f
C2337 VN.t16 AVSS 0.496456f
C2338 VN.n793 AVSS 0.239402f
C2339 VN.n794 AVSS 0.063168f
C2340 VN.n795 AVSS 0.035125f
C2341 VN.n796 AVSS 0.064726f
C2342 VN.n797 AVSS 0.064726f
C2343 VN.t56 AVSS 0.496456f
C2344 VN.n798 AVSS 0.239398f
C2345 VN.n799 AVSS 0.053679f
C2346 VN.n800 AVSS 0.035125f
C2347 VN.n801 AVSS 0.053679f
C2348 VN.n802 AVSS 0.053679f
C2349 VN.n803 AVSS 0.035125f
C2350 VN.n804 AVSS 0.073628f
C2351 VN.n805 AVSS 0.053679f
C2352 VN.n806 AVSS 0.188544f
C2353 VN.n807 AVSS 0.188544f
C2354 VN.n808 AVSS 0.082083f
C2355 VN.n809 AVSS 0.035125f
C2356 VN.n810 AVSS 0.064726f
C2357 VN.n811 AVSS 0.206949f
C2358 VN.n812 AVSS 0.227348f
C2359 VN.n813 AVSS 0.075617f
C2360 VN.n814 AVSS 0.035125f
C2361 VN.n815 AVSS 0.063168f
C2362 VN.n816 AVSS 0.063168f
C2363 VN.n817 AVSS 0.221877f
C2364 VN.n818 AVSS 0.074622f
C2365 VN.t41 AVSS 0.496456f
C2366 VN.n819 AVSS 0.239402f
C2367 VN.n820 AVSS 0.090542f
C2368 VN.n821 AVSS 0.39827f
C2369 VN.n822 AVSS 0.39827f
C2370 VN.n823 AVSS 0.089547f
C2371 VN.n824 AVSS 0.39827f
C2372 VN.n825 AVSS 0.035125f
C2373 VN.n826 AVSS 0.053679f
C2374 VN.n827 AVSS 0.188544f
C2375 VN.n828 AVSS 0.188544f
C2376 VN.n829 AVSS 0.082083f
C2377 VN.n830 AVSS 0.035125f
C2378 VN.n831 AVSS 0.064726f
C2379 VN.n832 AVSS 0.064726f
C2380 VN.n833 AVSS 0.227348f
C2381 VN.n834 AVSS 0.075617f
C2382 VN.t58 AVSS 0.496456f
C2383 VN.n835 AVSS 0.239402f
C2384 VN.n836 AVSS 0.207948f
C2385 VN.n837 AVSS 0.063168f
C2386 VN.n838 AVSS 0.063168f
C2387 VN.n839 AVSS 0.035125f
C2388 VN.n840 AVSS 0.074622f
C2389 VN.t81 AVSS 0.496456f
C2390 VN.n841 AVSS 0.239402f
C2391 VN.n842 AVSS 0.090542f
C2392 VN.n843 AVSS 0.282131f
C2393 VN.n844 AVSS 0.370227f
C2394 VN.n845 AVSS 7.09337f
C2395 VN.n846 AVSS 7.09129f
C2396 VN.n847 AVSS 0.370227f
C2397 VN.n848 AVSS 0.12322f
C2398 VN.n849 AVSS 0.053728f
C2399 a_n13990_n6451.n0 AVSS 0.969528f
C2400 a_n13990_n6451.n1 AVSS 0.842154f
C2401 a_n13990_n6451.n2 AVSS 0.923689f
C2402 a_n13990_n6451.n3 AVSS 0.630999f
C2403 a_n13990_n6451.n4 AVSS 0.937198f
C2404 a_n13990_n6451.n5 AVSS 0.937197f
C2405 a_n13990_n6451.n6 AVSS 0.497665f
C2406 a_n13990_n6451.n7 AVSS 0.842154f
C2407 a_n13990_n6451.n8 AVSS 0.923689f
C2408 a_n13990_n6451.n9 AVSS 1.10039f
C2409 a_n13990_n6451.n10 AVSS 0.969528f
C2410 a_n13990_n6451.n11 AVSS 0.842154f
C2411 a_n13990_n6451.n12 AVSS 0.923689f
C2412 a_n13990_n6451.n13 AVSS 0.630999f
C2413 a_n13990_n6451.n14 AVSS 0.937198f
C2414 a_n13990_n6451.n15 AVSS 0.937197f
C2415 a_n13990_n6451.n16 AVSS 0.497665f
C2416 a_n13990_n6451.n17 AVSS 0.842154f
C2417 a_n13990_n6451.n18 AVSS 0.923689f
C2418 a_n13990_n6451.n19 AVSS 1.10039f
C2419 a_n13990_n6451.n20 AVSS 0.556333f
C2420 a_n13990_n6451.n21 AVSS 0.888363f
C2421 a_n13990_n6451.n22 AVSS 1.47271f
C2422 a_n13990_n6451.n23 AVSS 0.952191f
C2423 a_n13990_n6451.n24 AVSS 0.825245f
C2424 a_n13990_n6451.n25 AVSS 1.46532f
C2425 a_n13990_n6451.t56 AVSS 0.429175f
C2426 a_n13990_n6451.t108 AVSS 0.076655f
C2427 a_n13990_n6451.t84 AVSS 0.076655f
C2428 a_n13990_n6451.n26 AVSS 0.331846f
C2429 a_n13990_n6451.n27 AVSS 1.09234f
C2430 a_n13990_n6451.t85 AVSS 0.325318f
C2431 a_n13990_n6451.n28 AVSS 0.924587f
C2432 a_n13990_n6451.t71 AVSS 0.076655f
C2433 a_n13990_n6451.t133 AVSS 0.076655f
C2434 a_n13990_n6451.n29 AVSS 0.331846f
C2435 a_n13990_n6451.n30 AVSS 0.497993f
C2436 a_n13990_n6451.n31 AVSS 3.12728f
C2437 a_n13990_n6451.n32 AVSS 3.94907f
C2438 a_n13990_n6451.t105 AVSS 0.188932f
C2439 a_n13990_n6451.t103 AVSS 0.230522f
C2440 a_n13990_n6451.n33 AVSS 1.2354f
C2441 a_n13990_n6451.t124 AVSS 0.076655f
C2442 a_n13990_n6451.t64 AVSS 0.076655f
C2443 a_n13990_n6451.n34 AVSS 0.179401f
C2444 a_n13990_n6451.t121 AVSS 0.076655f
C2445 a_n13990_n6451.t63 AVSS 0.076655f
C2446 a_n13990_n6451.n35 AVSS 0.228235f
C2447 a_n13990_n6451.n36 AVSS 0.519478f
C2448 a_n13990_n6451.n37 AVSS 1.13555f
C2449 a_n13990_n6451.t134 AVSS 0.43522f
C2450 a_n13990_n6451.t65 AVSS 0.076655f
C2451 a_n13990_n6451.t106 AVSS 0.076655f
C2452 a_n13990_n6451.n38 AVSS 0.331846f
C2453 a_n13990_n6451.n39 AVSS 0.974161f
C2454 a_n13990_n6451.n40 AVSS 0.746834f
C2455 a_n13990_n6451.t80 AVSS 0.188932f
C2456 a_n13990_n6451.t82 AVSS 0.230522f
C2457 a_n13990_n6451.n41 AVSS 1.2354f
C2458 a_n13990_n6451.t86 AVSS 0.076655f
C2459 a_n13990_n6451.t59 AVSS 0.076655f
C2460 a_n13990_n6451.n42 AVSS 0.179401f
C2461 a_n13990_n6451.t88 AVSS 0.076655f
C2462 a_n13990_n6451.t61 AVSS 0.076655f
C2463 a_n13990_n6451.n43 AVSS 0.228235f
C2464 a_n13990_n6451.n44 AVSS 0.519478f
C2465 a_n13990_n6451.n45 AVSS 1.13555f
C2466 a_n13990_n6451.t81 AVSS 0.429175f
C2467 a_n13990_n6451.t75 AVSS 0.076655f
C2468 a_n13990_n6451.t68 AVSS 0.076655f
C2469 a_n13990_n6451.n46 AVSS 0.331846f
C2470 a_n13990_n6451.n47 AVSS 1.09234f
C2471 a_n13990_n6451.t130 AVSS 0.325318f
C2472 a_n13990_n6451.n48 AVSS 0.924535f
C2473 a_n13990_n6451.t113 AVSS 0.322533f
C2474 a_n13990_n6451.n49 AVSS 0.837697f
C2475 a_n13990_n6451.t58 AVSS 0.322533f
C2476 a_n13990_n6451.n50 AVSS 0.837697f
C2477 a_n13990_n6451.t95 AVSS 0.325318f
C2478 a_n13990_n6451.n51 AVSS 0.924535f
C2479 a_n13990_n6451.t137 AVSS 0.076655f
C2480 a_n13990_n6451.t118 AVSS 0.076655f
C2481 a_n13990_n6451.n52 AVSS 0.331846f
C2482 a_n13990_n6451.n53 AVSS 0.630758f
C2483 a_n13990_n6451.t74 AVSS 0.322533f
C2484 a_n13990_n6451.n54 AVSS 0.93037f
C2485 a_n13990_n6451.t77 AVSS 0.325227f
C2486 a_n13990_n6451.n55 AVSS 0.937996f
C2487 a_n13990_n6451.t119 AVSS 0.076655f
C2488 a_n13990_n6451.t73 AVSS 0.076655f
C2489 a_n13990_n6451.n56 AVSS 0.331846f
C2490 a_n13990_n6451.n57 AVSS 0.497993f
C2491 a_n13990_n6451.n58 AVSS 0.746834f
C2492 a_n13990_n6451.n59 AVSS 4.40324f
C2493 a_n13990_n6451.n60 AVSS 1.45516f
C2494 a_n13990_n6451.t109 AVSS 0.188932f
C2495 a_n13990_n6451.t110 AVSS 0.230522f
C2496 a_n13990_n6451.n61 AVSS 0.675571f
C2497 a_n13990_n6451.n62 AVSS 1.38083f
C2498 a_n13990_n6451.t139 AVSS 0.076655f
C2499 a_n13990_n6451.t111 AVSS 0.076655f
C2500 a_n13990_n6451.n63 AVSS 0.179401f
C2501 a_n13990_n6451.t141 AVSS 0.076655f
C2502 a_n13990_n6451.t112 AVSS 0.076655f
C2503 a_n13990_n6451.n64 AVSS 0.228235f
C2504 a_n13990_n6451.n65 AVSS 0.519478f
C2505 a_n13990_n6451.n66 AVSS 0.902893f
C2506 a_n13990_n6451.n67 AVSS 4.88139f
C2507 a_n13990_n6451.t116 AVSS 0.433213f
C2508 a_n13990_n6451.t90 AVSS 0.076655f
C2509 a_n13990_n6451.t127 AVSS 0.076655f
C2510 a_n13990_n6451.n68 AVSS 0.331171f
C2511 a_n13990_n6451.t70 AVSS 0.324657f
C2512 a_n13990_n6451.t55 AVSS 0.324236f
C2513 a_n13990_n6451.n69 AVSS 0.213675f
C2514 a_n13990_n6451.t91 AVSS 0.076655f
C2515 a_n13990_n6451.t83 AVSS 0.076655f
C2516 a_n13990_n6451.n70 AVSS 0.331171f
C2517 a_n13990_n6451.t114 AVSS 0.324657f
C2518 a_n13990_n6451.t104 AVSS 0.324657f
C2519 a_n13990_n6451.t69 AVSS 0.076655f
C2520 a_n13990_n6451.t131 AVSS 0.076655f
C2521 a_n13990_n6451.n71 AVSS 0.331171f
C2522 a_n13990_n6451.t97 AVSS 0.324657f
C2523 a_n13990_n6451.t93 AVSS 0.324236f
C2524 a_n13990_n6451.t129 AVSS 0.076655f
C2525 a_n13990_n6451.t117 AVSS 0.076655f
C2526 a_n13990_n6451.n72 AVSS 0.331171f
C2527 a_n13990_n6451.t57 AVSS 0.433794f
C2528 a_n13990_n6451.n73 AVSS 0.213675f
C2529 a_n13990_n6451.n74 AVSS 3.12728f
C2530 a_n13990_n6451.t62 AVSS 0.325227f
C2531 a_n13990_n6451.n75 AVSS 0.937996f
C2532 a_n13990_n6451.t89 AVSS 0.322533f
C2533 a_n13990_n6451.n76 AVSS 0.93037f
C2534 a_n13990_n6451.t115 AVSS 0.076655f
C2535 a_n13990_n6451.t78 AVSS 0.076655f
C2536 a_n13990_n6451.n77 AVSS 0.331846f
C2537 a_n13990_n6451.n78 AVSS 0.630758f
C2538 a_n13990_n6451.t107 AVSS 0.325318f
C2539 a_n13990_n6451.n79 AVSS 0.924535f
C2540 a_n13990_n6451.t135 AVSS 0.322533f
C2541 a_n13990_n6451.n80 AVSS 0.837697f
C2542 a_n13990_n6451.t122 AVSS 0.43522f
C2543 a_n13990_n6451.t66 AVSS 0.076655f
C2544 a_n13990_n6451.t126 AVSS 0.076655f
C2545 a_n13990_n6451.n81 AVSS 0.331846f
C2546 a_n13990_n6451.n82 AVSS 0.974161f
C2547 a_n13990_n6451.n83 AVSS 0.213683f
C2548 a_n13990_n6451.n84 AVSS 2.81125f
C2549 a_n13990_n6451.n85 AVSS 5.37523f
C2550 a_n13990_n6451.t26 AVSS 0.073005f
C2551 a_n13990_n6451.t6 AVSS 0.073005f
C2552 a_n13990_n6451.n86 AVSS 0.373178f
C2553 a_n13990_n6451.n87 AVSS 1.61957f
C2554 a_n13990_n6451.t4 AVSS 0.188802f
C2555 a_n13990_n6451.t11 AVSS 0.227347f
C2556 a_n13990_n6451.n88 AVSS 1.13041f
C2557 a_n13990_n6451.t24 AVSS 0.073005f
C2558 a_n13990_n6451.t49 AVSS 0.073005f
C2559 a_n13990_n6451.n89 AVSS 0.168553f
C2560 a_n13990_n6451.t17 AVSS 0.073005f
C2561 a_n13990_n6451.t12 AVSS 0.073005f
C2562 a_n13990_n6451.n90 AVSS 0.212607f
C2563 a_n13990_n6451.n91 AVSS 0.533434f
C2564 a_n13990_n6451.n92 AVSS 1.04553f
C2565 a_n13990_n6451.t10 AVSS 0.431942f
C2566 a_n13990_n6451.t25 AVSS 0.073005f
C2567 a_n13990_n6451.t22 AVSS 0.073005f
C2568 a_n13990_n6451.n93 AVSS 0.309391f
C2569 a_n13990_n6451.t8 AVSS 0.317687f
C2570 a_n13990_n6451.n94 AVSS 0.949857f
C2571 a_n13990_n6451.t30 AVSS 0.073005f
C2572 a_n13990_n6451.t21 AVSS 0.073005f
C2573 a_n13990_n6451.n95 AVSS 0.309391f
C2574 a_n13990_n6451.t7 AVSS 0.073005f
C2575 a_n13990_n6451.t28 AVSS 0.073005f
C2576 a_n13990_n6451.n96 AVSS 0.309391f
C2577 a_n13990_n6451.t5 AVSS 0.317687f
C2578 a_n13990_n6451.n97 AVSS 0.949857f
C2579 a_n13990_n6451.t51 AVSS 0.317687f
C2580 a_n13990_n6451.n98 AVSS 1.03306f
C2581 a_n13990_n6451.n99 AVSS 1.04012f
C2582 a_n13990_n6451.n100 AVSS 4.74525f
C2583 a_n13990_n6451.n101 AVSS 1.23914f
C2584 a_n13990_n6451.t20 AVSS 0.188802f
C2585 a_n13990_n6451.t18 AVSS 0.227347f
C2586 a_n13990_n6451.n102 AVSS 0.651755f
C2587 a_n13990_n6451.n103 AVSS 1.16321f
C2588 a_n13990_n6451.t13 AVSS 0.073005f
C2589 a_n13990_n6451.t9 AVSS 0.073005f
C2590 a_n13990_n6451.n104 AVSS 0.168553f
C2591 a_n13990_n6451.t53 AVSS 0.073005f
C2592 a_n13990_n6451.t3 AVSS 0.073005f
C2593 a_n13990_n6451.n105 AVSS 0.212607f
C2594 a_n13990_n6451.n106 AVSS 0.533434f
C2595 a_n13990_n6451.n107 AVSS 0.846593f
C2596 a_n13990_n6451.n108 AVSS 5.16107f
C2597 a_n13990_n6451.t29 AVSS 0.073005f
C2598 a_n13990_n6451.t52 AVSS 0.073005f
C2599 a_n13990_n6451.n109 AVSS 0.47617f
C2600 a_n13990_n6451.t50 AVSS 0.316937f
C2601 a_n13990_n6451.n110 AVSS 1.5065f
C2602 a_n13990_n6451.t1 AVSS 0.314232f
C2603 a_n13990_n6451.n111 AVSS 0.831997f
C2604 a_n13990_n6451.n112 AVSS 0.210773f
C2605 a_n13990_n6451.t19 AVSS 0.073005f
C2606 a_n13990_n6451.t2 AVSS 0.073005f
C2607 a_n13990_n6451.n113 AVSS 0.309971f
C2608 a_n13990_n6451.n114 AVSS 0.927634f
C2609 a_n13990_n6451.t14 AVSS 0.073005f
C2610 a_n13990_n6451.t0 AVSS 0.073005f
C2611 a_n13990_n6451.n115 AVSS 0.309971f
C2612 a_n13990_n6451.n116 AVSS 1.05597f
C2613 a_n13990_n6451.t27 AVSS 0.316937f
C2614 a_n13990_n6451.n117 AVSS 0.92047f
C2615 a_n13990_n6451.t15 AVSS 0.314232f
C2616 a_n13990_n6451.n118 AVSS 0.831997f
C2617 a_n13990_n6451.t23 AVSS 0.073005f
C2618 a_n13990_n6451.t16 AVSS 0.073005f
C2619 a_n13990_n6451.n119 AVSS 0.373767f
C2620 a_n13990_n6451.n120 AVSS 0.790666f
C2621 a_n13990_n6451.n121 AVSS 4.36492f
C2622 a_n13990_n6451.n122 AVSS 5.60327f
C2623 a_n13990_n6451.t47 AVSS 0.073005f
C2624 a_n13990_n6451.t34 AVSS 0.073005f
C2625 a_n13990_n6451.n123 AVSS 0.426576f
C2626 a_n13990_n6451.t46 AVSS 0.275089f
C2627 a_n13990_n6451.t42 AVSS 0.073005f
C2628 a_n13990_n6451.t48 AVSS 0.073005f
C2629 a_n13990_n6451.n124 AVSS 0.261791f
C2630 a_n13990_n6451.t41 AVSS 0.275089f
C2631 a_n13990_n6451.n125 AVSS 3.22126f
C2632 a_n13990_n6451.t45 AVSS 0.073005f
C2633 a_n13990_n6451.t33 AVSS 0.073005f
C2634 a_n13990_n6451.n126 AVSS 0.197177f
C2635 a_n13990_n6451.t39 AVSS 0.073005f
C2636 a_n13990_n6451.t43 AVSS 0.073005f
C2637 a_n13990_n6451.n127 AVSS 0.180875f
C2638 a_n13990_n6451.n128 AVSS 1.11951f
C2639 a_n13990_n6451.t44 AVSS 0.213949f
C2640 a_n13990_n6451.t38 AVSS 0.199722f
C2641 a_n13990_n6451.n129 AVSS 0.664361f
C2642 a_n13990_n6451.n130 AVSS 1.44653f
C2643 a_n13990_n6451.n131 AVSS 2.99913f
C2644 a_n13990_n6451.t36 AVSS 0.381078f
C2645 a_n13990_n6451.t40 AVSS 0.073005f
C2646 a_n13990_n6451.t35 AVSS 0.073005f
C2647 a_n13990_n6451.n132 AVSS 0.262553f
C2648 a_n13990_n6451.n133 AVSS 1.43556f
C2649 a_n13990_n6451.t32 AVSS 0.073005f
C2650 a_n13990_n6451.t37 AVSS 0.073005f
C2651 a_n13990_n6451.n134 AVSS 0.262553f
C2652 a_n13990_n6451.n135 AVSS 0.991537f
C2653 a_n13990_n6451.t31 AVSS 0.275734f
C2654 a_n13990_n6451.n136 AVSS 0.554014f
C2655 a_n13990_n6451.n137 AVSS 8.83141f
C2656 a_n13990_n6451.n138 AVSS 12.0991f
C2657 a_n13990_n6451.t72 AVSS 0.433213f
C2658 a_n13990_n6451.t128 AVSS 0.076655f
C2659 a_n13990_n6451.t100 AVSS 0.076655f
C2660 a_n13990_n6451.n139 AVSS 0.331171f
C2661 a_n13990_n6451.t101 AVSS 0.324657f
C2662 a_n13990_n6451.t67 AVSS 0.324236f
C2663 a_n13990_n6451.n140 AVSS 0.213675f
C2664 a_n13990_n6451.t87 AVSS 0.076655f
C2665 a_n13990_n6451.t54 AVSS 0.076655f
C2666 a_n13990_n6451.n141 AVSS 0.331171f
C2667 a_n13990_n6451.t76 AVSS 0.324657f
C2668 a_n13990_n6451.t102 AVSS 0.324657f
C2669 a_n13990_n6451.t132 AVSS 0.076655f
C2670 a_n13990_n6451.t92 AVSS 0.076655f
C2671 a_n13990_n6451.n142 AVSS 0.331171f
C2672 a_n13990_n6451.t120 AVSS 0.324657f
C2673 a_n13990_n6451.t60 AVSS 0.324236f
C2674 a_n13990_n6451.t79 AVSS 0.076655f
C2675 a_n13990_n6451.t138 AVSS 0.076655f
C2676 a_n13990_n6451.n143 AVSS 0.331171f
C2677 a_n13990_n6451.t136 AVSS 0.433794f
C2678 a_n13990_n6451.n144 AVSS 0.213675f
C2679 a_n13990_n6451.n145 AVSS 7.5285f
C2680 a_n13990_n6451.n146 AVSS 3.62772f
C2681 a_n13990_n6451.t96 AVSS 0.076655f
C2682 a_n13990_n6451.t125 AVSS 0.076655f
C2683 a_n13990_n6451.n147 AVSS 0.179401f
C2684 a_n13990_n6451.t94 AVSS 0.076655f
C2685 a_n13990_n6451.t123 AVSS 0.076655f
C2686 a_n13990_n6451.n148 AVSS 0.228235f
C2687 a_n13990_n6451.n149 AVSS 0.519478f
C2688 a_n13990_n6451.n150 AVSS 0.902893f
C2689 a_n13990_n6451.t99 AVSS 0.188932f
C2690 a_n13990_n6451.t98 AVSS 0.230522f
C2691 a_n13990_n6451.n151 AVSS 0.675571f
C2692 a_n13990_n6451.n152 AVSS 1.38083f
C2693 a_n13990_n6451.n153 AVSS 1.45516f
C2694 a_n13990_n6451.n154 AVSS 3.14957f
C2695 a_n13990_n6451.n155 AVSS 2.81125f
C2696 a_n13990_n6451.n156 AVSS 0.213644f
C2697 a_n13990_n6451.n157 AVSS 0.837684f
C2698 a_n13990_n6451.t140 AVSS 0.322533f
C2699 VP.t18 AVSS 0.643351f
C2700 VP.n0 AVSS 0.494836f
C2701 VP.n1 AVSS 0.022318f
C2702 VP.n2 AVSS 0.376256f
C2703 VP.n3 AVSS 4.56964f
C2704 VP.n4 AVSS 1.72503f
C2705 VP.n5 AVSS 0.376256f
C2706 VP.n6 AVSS 0.045518f
C2707 VP.n7 AVSS 0.077417f
C2708 VP.n8 AVSS 0.045518f
C2709 VP.n9 AVSS 0.07672f
C2710 VP.t51 AVSS 0.643351f
C2711 VP.n10 AVSS 0.335386f
C2712 VP.t25 AVSS 0.657177f
C2713 VP.n11 AVSS 0.479785f
C2714 VP.n12 AVSS 0.295681f
C2715 VP.n13 AVSS 0.081492f
C2716 VP.n14 AVSS 0.077417f
C2717 VP.n15 AVSS 0.022318f
C2718 VP.t14 AVSS 0.643351f
C2719 VP.n16 AVSS 0.251918f
C2720 VP.n17 AVSS 0.07672f
C2721 VP.n18 AVSS 0.081492f
C2722 VP.n19 AVSS 0.081492f
C2723 VP.n20 AVSS 0.045518f
C2724 VP.n21 AVSS 0.022318f
C2725 VP.t71 AVSS 0.643351f
C2726 VP.n22 AVSS 0.251918f
C2727 VP.n23 AVSS 0.215658f
C2728 VP.t59 AVSS 0.643351f
C2729 VP.n24 AVSS 0.520988f
C2730 VP.t53 AVSS 0.643351f
C2731 VP.n25 AVSS 0.428373f
C2732 VP.t80 AVSS 0.643351f
C2733 VP.n26 AVSS 0.519478f
C2734 VP.n27 AVSS 0.077417f
C2735 VP.n28 AVSS 0.081492f
C2736 VP.n29 AVSS 0.022318f
C2737 VP.n30 AVSS 0.081492f
C2738 VP.t58 AVSS 0.643351f
C2739 VP.n31 AVSS 0.251918f
C2740 VP.t27 AVSS 0.643351f
C2741 VP.n32 AVSS 0.285723f
C2742 VP.n33 AVSS 0.096423f
C2743 VP.n34 AVSS 0.022318f
C2744 VP.n35 AVSS 0.081492f
C2745 VP.t72 AVSS 0.643351f
C2746 VP.n36 AVSS 0.251918f
C2747 VP.t10 AVSS 0.643351f
C2748 VP.n37 AVSS 0.251918f
C2749 VP.n38 AVSS 0.081492f
C2750 VP.t44 AVSS 0.643351f
C2751 VP.n39 AVSS 0.251918f
C2752 VP.n40 AVSS 0.379927f
C2753 VP.n41 AVSS 0.045518f
C2754 VP.n42 AVSS 0.066083f
C2755 VP.n43 AVSS 0.045518f
C2756 VP.n44 AVSS 0.079684f
C2757 VP.n45 AVSS 0.081859f
C2758 VP.n46 AVSS 0.026154f
C2759 VP.n47 AVSS 0.045518f
C2760 VP.n48 AVSS 0.066083f
C2761 VP.n49 AVSS 0.083878f
C2762 VP.n50 AVSS 0.026503f
C2763 VP.n51 AVSS 0.081859f
C2764 VP.t28 AVSS 0.643351f
C2765 VP.n52 AVSS 0.251918f
C2766 VP.t11 AVSS 0.643351f
C2767 VP.n53 AVSS 0.251918f
C2768 VP.n54 AVSS 0.069562f
C2769 VP.n55 AVSS 0.02877f
C2770 VP.n56 AVSS 0.083878f
C2771 VP.t66 AVSS 0.643351f
C2772 VP.n57 AVSS 0.318134f
C2773 VP.t60 AVSS 0.652717f
C2774 VP.n58 AVSS 0.449407f
C2775 VP.n59 AVSS 0.251521f
C2776 VP.n60 AVSS 0.026503f
C2777 VP.n61 AVSS 0.079684f
C2778 VP.t73 AVSS 0.643351f
C2779 VP.n62 AVSS 0.251918f
C2780 VP.n63 AVSS 0.072535f
C2781 VP.n64 AVSS 0.083878f
C2782 VP.n65 AVSS 0.045518f
C2783 VP.n66 AVSS 0.069562f
C2784 VP.n67 AVSS 0.066083f
C2785 VP.n68 AVSS 0.066083f
C2786 VP.n69 AVSS 0.025806f
C2787 VP.n70 AVSS 0.045518f
C2788 VP.n71 AVSS 0.379927f
C2789 VP.n72 AVSS 0.215377f
C2790 VP.t61 AVSS 0.643351f
C2791 VP.n73 AVSS 0.524756f
C2792 VP.t55 AVSS 0.643351f
C2793 VP.n74 AVSS 0.428373f
C2794 VP.t82 AVSS 0.643351f
C2795 VP.n75 AVSS 0.525183f
C2796 VP.n76 AVSS 0.215299f
C2797 VP.n77 AVSS 0.145363f
C2798 VP.n78 AVSS 0.045518f
C2799 VP.n79 AVSS 0.026154f
C2800 VP.n80 AVSS 0.077766f
C2801 VP.t22 AVSS 0.643351f
C2802 VP.n81 AVSS 0.251918f
C2803 VP.n82 AVSS 0.072884f
C2804 VP.n83 AVSS 0.081859f
C2805 VP.n84 AVSS 0.045518f
C2806 VP.n85 AVSS 0.083878f
C2807 VP.n86 AVSS 0.079684f
C2808 VP.n87 AVSS 0.072535f
C2809 VP.t68 AVSS 0.643351f
C2810 VP.n88 AVSS 0.251918f
C2811 VP.n89 AVSS 0.02877f
C2812 VP.n90 AVSS 0.045518f
C2813 VP.n91 AVSS 0.069562f
C2814 VP.n92 AVSS 0.069562f
C2815 VP.n93 AVSS 0.066083f
C2816 VP.n94 AVSS 0.025806f
C2817 VP.t64 AVSS 0.643351f
C2818 VP.n95 AVSS 0.289294f
C2819 VP.n96 AVSS 0.517097f
C2820 VP.t67 AVSS 0.643351f
C2821 VP.n97 AVSS 0.282854f
C2822 VP.n98 AVSS 0.516911f
C2823 VP.n99 AVSS 0.045518f
C2824 VP.n100 AVSS 0.081859f
C2825 VP.n101 AVSS 0.077766f
C2826 VP.n102 AVSS 0.072884f
C2827 VP.t4 AVSS 0.643351f
C2828 VP.n103 AVSS 0.251918f
C2829 VP.n104 AVSS 0.026503f
C2830 VP.n105 AVSS 0.045518f
C2831 VP.n106 AVSS 0.083878f
C2832 VP.n107 AVSS 0.083878f
C2833 VP.n108 AVSS 0.072535f
C2834 VP.t23 AVSS 0.643351f
C2835 VP.n109 AVSS 0.251918f
C2836 VP.n110 AVSS 0.02877f
C2837 VP.n111 AVSS 0.066083f
C2838 VP.n112 AVSS 0.069562f
C2839 VP.n113 AVSS 0.069562f
C2840 VP.n114 AVSS 0.045518f
C2841 VP.n115 AVSS 0.025806f
C2842 VP.t46 AVSS 0.643351f
C2843 VP.n116 AVSS 0.251918f
C2844 VP.n117 AVSS 0.215377f
C2845 VP.t32 AVSS 0.643351f
C2846 VP.n118 AVSS 0.524756f
C2847 VP.t2 AVSS 0.643351f
C2848 VP.n119 AVSS 0.428373f
C2849 VP.t30 AVSS 0.643351f
C2850 VP.n120 AVSS 0.525183f
C2851 VP.n121 AVSS 0.072884f
C2852 VP.n122 AVSS 0.083878f
C2853 VP.t76 AVSS 0.643351f
C2854 VP.n123 AVSS 0.251918f
C2855 VP.t35 AVSS 0.643351f
C2856 VP.n124 AVSS 0.323197f
C2857 VP.t7 AVSS 0.656201f
C2858 VP.n125 AVSS 0.479343f
C2859 VP.n126 AVSS 0.293659f
C2860 VP.n127 AVSS 0.072535f
C2861 VP.n128 AVSS 0.079684f
C2862 VP.n129 AVSS 0.026503f
C2863 VP.n130 AVSS 0.045518f
C2864 VP.n131 AVSS 0.081859f
C2865 VP.n132 AVSS 0.081859f
C2866 VP.n133 AVSS 0.077766f
C2867 VP.n134 AVSS 0.026154f
C2868 VP.t83 AVSS 0.643351f
C2869 VP.n135 AVSS 0.251918f
C2870 VP.n136 AVSS 0.215299f
C2871 VP.n137 AVSS 0.145363f
C2872 VP.n138 AVSS 1.72503f
C2873 VP.n139 AVSS 6.87741f
C2874 VP.n140 AVSS 0.470596f
C2875 VP.n141 AVSS 0.022318f
C2876 VP.n142 AVSS 0.081492f
C2877 VP.t48 AVSS 0.643351f
C2878 VP.n143 AVSS 0.251918f
C2879 VP.t12 AVSS 0.643351f
C2880 VP.n144 AVSS 0.251918f
C2881 VP.n145 AVSS 0.081492f
C2882 VP.t24 AVSS 0.643351f
C2883 VP.n146 AVSS 0.315255f
C2884 VP.t84 AVSS 0.652002f
C2885 VP.n147 AVSS 0.454236f
C2886 VP.n148 AVSS 0.249774f
C2887 VP.n149 AVSS 0.022318f
C2888 VP.n150 AVSS 0.077417f
C2889 VP.n151 AVSS 0.07672f
C2890 VP.n152 AVSS 0.081492f
C2891 VP.n153 AVSS 0.045518f
C2892 VP.n154 AVSS 0.022318f
C2893 VP.n155 AVSS 0.077417f
C2894 VP.n156 AVSS 0.07672f
C2895 VP.n157 AVSS 0.081492f
C2896 VP.n158 AVSS 0.045518f
C2897 VP.n159 AVSS 0.139857f
C2898 VP.n160 AVSS 0.215076f
C2899 VP.t29 AVSS 0.643351f
C2900 VP.n161 AVSS 0.519478f
C2901 VP.t0 AVSS 0.643351f
C2902 VP.n162 AVSS 0.428373f
C2903 VP.t31 AVSS 0.643351f
C2904 VP.n163 AVSS 0.520988f
C2905 VP.n164 AVSS 0.215658f
C2906 VP.n165 AVSS 0.376256f
C2907 VP.n166 AVSS 0.045518f
C2908 VP.n167 AVSS 0.022318f
C2909 VP.n168 AVSS 0.077417f
C2910 VP.n169 AVSS 0.07672f
C2911 VP.n170 AVSS 0.081492f
C2912 VP.n171 AVSS 0.045518f
C2913 VP.n172 AVSS 0.022318f
C2914 VP.n173 AVSS 0.077417f
C2915 VP.n174 AVSS 0.07672f
C2916 VP.n175 AVSS 0.081492f
C2917 VP.n176 AVSS 0.045518f
C2918 VP.n177 AVSS 0.081492f
C2919 VP.n178 AVSS 0.077417f
C2920 VP.n179 AVSS 0.07672f
C2921 VP.t37 AVSS 0.643351f
C2922 VP.n180 AVSS 0.309237f
C2923 VP.n181 AVSS 0.527032f
C2924 VP.n182 AVSS 0.519762f
C2925 VP.n183 AVSS 0.045518f
C2926 VP.n184 AVSS 0.022318f
C2927 VP.n185 AVSS 0.077417f
C2928 VP.n186 AVSS 0.07672f
C2929 VP.n187 AVSS 0.081492f
C2930 VP.n188 AVSS 0.045518f
C2931 VP.n189 AVSS 0.081492f
C2932 VP.n190 AVSS 0.077417f
C2933 VP.n191 AVSS 0.07672f
C2934 VP.t50 AVSS 0.643351f
C2935 VP.n192 AVSS 0.251918f
C2936 VP.n193 AVSS 0.022318f
C2937 VP.n194 AVSS 0.045518f
C2938 VP.n195 AVSS 0.081492f
C2939 VP.n196 AVSS 0.081492f
C2940 VP.n197 AVSS 0.07672f
C2941 VP.t86 AVSS 0.643351f
C2942 VP.n198 AVSS 0.251918f
C2943 VP.n199 AVSS 0.022318f
C2944 VP.n200 AVSS 0.215076f
C2945 VP.n201 AVSS 0.139857f
C2946 VP.n202 AVSS 0.470596f
C2947 VP.n203 AVSS 6.87741f
C2948 VP.n204 AVSS 0.379927f
C2949 VP.n205 AVSS 0.045518f
C2950 VP.n206 AVSS 0.066083f
C2951 VP.n207 AVSS 0.045518f
C2952 VP.n208 AVSS 0.079684f
C2953 VP.t85 AVSS 0.652717f
C2954 VP.n209 AVSS 0.449407f
C2955 VP.t33 AVSS 0.643351f
C2956 VP.n210 AVSS 0.318134f
C2957 VP.n211 AVSS 0.026503f
C2958 VP.n212 AVSS 0.251521f
C2959 VP.n213 AVSS 0.083878f
C2960 VP.n214 AVSS 0.083878f
C2961 VP.n215 AVSS 0.072535f
C2962 VP.t57 AVSS 0.643351f
C2963 VP.n216 AVSS 0.251918f
C2964 VP.n217 AVSS 0.02877f
C2965 VP.n218 AVSS 0.066083f
C2966 VP.n219 AVSS 0.069562f
C2967 VP.n220 AVSS 0.069562f
C2968 VP.n221 AVSS 0.045518f
C2969 VP.n222 AVSS 0.025806f
C2970 VP.t56 AVSS 0.643351f
C2971 VP.n223 AVSS 0.251918f
C2972 VP.n224 AVSS 0.215377f
C2973 VP.t36 AVSS 0.643351f
C2974 VP.n225 AVSS 0.524756f
C2975 VP.t17 AVSS 0.643351f
C2976 VP.n226 AVSS 0.428373f
C2977 VP.t77 AVSS 0.643351f
C2978 VP.n227 AVSS 0.525183f
C2979 VP.n228 AVSS 0.072884f
C2980 VP.n229 AVSS 0.083878f
C2981 VP.t70 AVSS 0.643351f
C2982 VP.n230 AVSS 0.251918f
C2983 VP.t8 AVSS 0.643351f
C2984 VP.n231 AVSS 0.251918f
C2985 VP.n232 AVSS 0.069562f
C2986 VP.n233 AVSS 0.025806f
C2987 VP.n234 AVSS 0.045518f
C2988 VP.n235 AVSS 0.072884f
C2989 VP.n236 AVSS 0.083878f
C2990 VP.t26 AVSS 0.643351f
C2991 VP.n237 AVSS 0.251918f
C2992 VP.t63 AVSS 0.643351f
C2993 VP.n238 AVSS 0.251918f
C2994 VP.n239 AVSS 0.069562f
C2995 VP.n240 AVSS 0.025806f
C2996 VP.n241 AVSS 0.479772f
C2997 VP.t34 AVSS 0.643351f
C2998 VP.n242 AVSS 0.251918f
C2999 VP.t6 AVSS 0.643351f
C3000 VP.n243 AVSS 0.251918f
C3001 VP.n244 AVSS 0.081859f
C3002 VP.t75 AVSS 0.643351f
C3003 VP.n245 AVSS 0.251918f
C3004 VP.n246 AVSS 0.083878f
C3005 VP.t15 AVSS 0.643351f
C3006 VP.n247 AVSS 0.323197f
C3007 VP.t19 AVSS 0.656201f
C3008 VP.n248 AVSS 0.479343f
C3009 VP.n249 AVSS 0.293659f
C3010 VP.n250 AVSS 0.072535f
C3011 VP.n251 AVSS 0.079684f
C3012 VP.n252 AVSS 0.026503f
C3013 VP.n253 AVSS 0.045518f
C3014 VP.n254 AVSS 0.081859f
C3015 VP.n255 AVSS 0.072884f
C3016 VP.n256 AVSS 0.077766f
C3017 VP.n257 AVSS 0.026154f
C3018 VP.n258 AVSS 0.045518f
C3019 VP.n259 AVSS 0.145363f
C3020 VP.n260 AVSS 0.215299f
C3021 VP.t16 AVSS 0.643351f
C3022 VP.n261 AVSS 0.525183f
C3023 VP.t45 AVSS 0.643351f
C3024 VP.n262 AVSS 0.428373f
C3025 VP.t42 AVSS 0.643351f
C3026 VP.n263 AVSS 0.524756f
C3027 VP.n264 AVSS 0.215377f
C3028 VP.n265 AVSS 0.379927f
C3029 VP.n266 AVSS 0.045518f
C3030 VP.n267 AVSS 0.069562f
C3031 VP.n268 AVSS 0.066083f
C3032 VP.n269 AVSS 0.066083f
C3033 VP.n270 AVSS 0.02877f
C3034 VP.n271 AVSS 0.045518f
C3035 VP.n272 AVSS 0.083878f
C3036 VP.n273 AVSS 0.072535f
C3037 VP.n274 AVSS 0.079684f
C3038 VP.n275 AVSS 0.026503f
C3039 VP.n276 AVSS 0.045518f
C3040 VP.n277 AVSS 0.081859f
C3041 VP.n278 AVSS 0.081859f
C3042 VP.n279 AVSS 0.077766f
C3043 VP.n280 AVSS 0.026154f
C3044 VP.t52 AVSS 0.643351f
C3045 VP.n281 AVSS 0.282854f
C3046 VP.n282 AVSS 0.516911f
C3047 VP.t79 AVSS 0.643351f
C3048 VP.n283 AVSS 0.289294f
C3049 VP.n284 AVSS 0.517097f
C3050 VP.n285 AVSS 0.045518f
C3051 VP.n286 AVSS 0.069562f
C3052 VP.n287 AVSS 0.066083f
C3053 VP.n288 AVSS 0.066083f
C3054 VP.n289 AVSS 0.02877f
C3055 VP.n290 AVSS 0.045518f
C3056 VP.n291 AVSS 0.083878f
C3057 VP.n292 AVSS 0.072535f
C3058 VP.n293 AVSS 0.079684f
C3059 VP.n294 AVSS 0.026503f
C3060 VP.n295 AVSS 0.045518f
C3061 VP.n296 AVSS 0.081859f
C3062 VP.n297 AVSS 0.081859f
C3063 VP.n298 AVSS 0.077766f
C3064 VP.n299 AVSS 0.026154f
C3065 VP.t1 AVSS 0.643351f
C3066 VP.n300 AVSS 0.251918f
C3067 VP.n301 AVSS 0.215299f
C3068 VP.n302 AVSS 0.145363f
C3069 VP.n303 AVSS 0.479772f
C3070 VP.n304 AVSS 4.56964f
C3071 VP.n305 AVSS 0.376256f
C3072 VP.n306 AVSS 0.045518f
C3073 VP.n307 AVSS 0.077417f
C3074 VP.n308 AVSS 0.045518f
C3075 VP.n309 AVSS 0.07672f
C3076 VP.t13 AVSS 0.643351f
C3077 VP.n310 AVSS 0.335386f
C3078 VP.t69 AVSS 0.657177f
C3079 VP.n311 AVSS 0.479785f
C3080 VP.n312 AVSS 0.295681f
C3081 VP.n313 AVSS 0.081492f
C3082 VP.n314 AVSS 0.077417f
C3083 VP.n315 AVSS 0.022318f
C3084 VP.t41 AVSS 0.643351f
C3085 VP.n316 AVSS 0.251918f
C3086 VP.n317 AVSS 0.07672f
C3087 VP.n318 AVSS 0.081492f
C3088 VP.n319 AVSS 0.081492f
C3089 VP.n320 AVSS 0.045518f
C3090 VP.n321 AVSS 0.022318f
C3091 VP.t40 AVSS 0.643351f
C3092 VP.n322 AVSS 0.251918f
C3093 VP.n323 AVSS 0.215658f
C3094 VP.t38 AVSS 0.643351f
C3095 VP.n324 AVSS 0.520988f
C3096 VP.t20 AVSS 0.643351f
C3097 VP.n325 AVSS 0.428373f
C3098 VP.t78 AVSS 0.643351f
C3099 VP.n326 AVSS 0.519478f
C3100 VP.n327 AVSS 0.077417f
C3101 VP.n328 AVSS 0.081492f
C3102 VP.n329 AVSS 0.022318f
C3103 VP.n330 AVSS 0.081492f
C3104 VP.t87 AVSS 0.643351f
C3105 VP.n331 AVSS 0.251918f
C3106 VP.t65 AVSS 0.643351f
C3107 VP.n332 AVSS 0.285723f
C3108 VP.n333 AVSS 0.096423f
C3109 VP.n334 AVSS 0.022318f
C3110 VP.n335 AVSS 0.081492f
C3111 VP.t9 AVSS 0.643351f
C3112 VP.n336 AVSS 0.251918f
C3113 VP.t49 AVSS 0.643351f
C3114 VP.n337 AVSS 0.251918f
C3115 VP.n338 AVSS 0.081492f
C3116 VP.t47 AVSS 0.643351f
C3117 VP.n339 AVSS 0.428373f
C3118 VP.t43 AVSS 0.643351f
C3119 VP.n340 AVSS 0.520988f
C3120 VP.n341 AVSS 0.215658f
C3121 VP.t21 AVSS 0.643351f
C3122 VP.n342 AVSS 0.251918f
C3123 VP.n343 AVSS 0.045518f
C3124 VP.n344 AVSS 0.022318f
C3125 VP.n345 AVSS 0.077417f
C3126 VP.n346 AVSS 0.07672f
C3127 VP.n347 AVSS 0.081492f
C3128 VP.n348 AVSS 0.045518f
C3129 VP.n349 AVSS 0.022318f
C3130 VP.n350 AVSS 0.077417f
C3131 VP.n351 AVSS 0.07672f
C3132 VP.n352 AVSS 0.081492f
C3133 VP.n353 AVSS 0.045518f
C3134 VP.n354 AVSS 0.081492f
C3135 VP.n355 AVSS 0.077417f
C3136 VP.n356 AVSS 0.07672f
C3137 VP.t39 AVSS 0.643351f
C3138 VP.n357 AVSS 0.309237f
C3139 VP.n358 AVSS 0.527032f
C3140 VP.n359 AVSS 0.519762f
C3141 VP.n360 AVSS 0.045518f
C3142 VP.n361 AVSS 0.022318f
C3143 VP.n362 AVSS 0.077417f
C3144 VP.n363 AVSS 0.07672f
C3145 VP.n364 AVSS 0.081492f
C3146 VP.n365 AVSS 0.045518f
C3147 VP.n366 AVSS 0.081492f
C3148 VP.n367 AVSS 0.077417f
C3149 VP.n368 AVSS 0.07672f
C3150 VP.t54 AVSS 0.643351f
C3151 VP.n369 AVSS 0.251918f
C3152 VP.n370 AVSS 0.022318f
C3153 VP.n371 AVSS 0.045518f
C3154 VP.n372 AVSS 0.081492f
C3155 VP.n373 AVSS 0.081492f
C3156 VP.n374 AVSS 0.07672f
C3157 VP.t74 AVSS 0.643351f
C3158 VP.n375 AVSS 0.251918f
C3159 VP.n376 AVSS 0.022318f
C3160 VP.n377 AVSS 0.215076f
C3161 VP.n378 AVSS 0.139857f
C3162 VP.n379 AVSS 0.470596f
C3163 VP.n380 AVSS 8.79061f
C3164 VP.n381 AVSS 8.714661f
C3165 VP.n382 AVSS 0.470596f
C3166 VP.n383 AVSS 0.081492f
C3167 VP.t81 AVSS 0.643351f
C3168 VP.n384 AVSS 0.251918f
C3169 VP.t62 AVSS 0.643351f
C3170 VP.n385 AVSS 0.251918f
C3171 VP.n386 AVSS 0.081492f
C3172 VP.t3 AVSS 0.643351f
C3173 VP.n387 AVSS 0.315255f
C3174 VP.t5 AVSS 0.652002f
C3175 VP.n388 AVSS 0.454235f
C3176 VP.n389 AVSS 0.249774f
C3177 VP.n390 AVSS 0.022318f
C3178 VP.n391 AVSS 0.077417f
C3179 VP.n392 AVSS 0.07672f
C3180 VP.n393 AVSS 0.081492f
C3181 VP.n394 AVSS 0.045518f
C3182 VP.n395 AVSS 0.022318f
C3183 VP.n396 AVSS 0.077417f
C3184 VP.n397 AVSS 0.07672f
C3185 VP.n398 AVSS 0.081492f
C3186 VP.n399 AVSS 0.045518f
C3187 VP.n400 AVSS 0.139857f
C3188 VP.n401 AVSS 0.044114f
C3189 a_n11317_n20927.t1 AVSS 0.227029p
C3190 a_n11317_n20927.t3 AVSS 0.587411f
C3191 a_n11317_n20927.t0 AVSS 2.58643f
C3192 a_n11317_n20927.t5 AVSS 0.339324f
C3193 a_n11317_n20927.t4 AVSS 3.45836f
C3194 a_n13990_8177.n0 AVSS 1.70465f
C3195 a_n13990_8177.n1 AVSS 1.49104f
C3196 a_n13990_8177.n2 AVSS 0.962831f
C3197 a_n13990_8177.n3 AVSS 1.70465f
C3198 a_n13990_8177.n4 AVSS 1.49104f
C3199 a_n13990_8177.n5 AVSS 0.962831f
C3200 a_n13990_8177.n6 AVSS 1.77854f
C3201 a_n13990_8177.n7 AVSS 1.25797f
C3202 a_n13990_8177.n8 AVSS 1.19957f
C3203 a_n13990_8177.n9 AVSS 1.77854f
C3204 a_n13990_8177.n10 AVSS 1.25797f
C3205 a_n13990_8177.n11 AVSS 0.91508f
C3206 a_n13990_8177.n12 AVSS 0.833972f
C3207 a_n13990_8177.n13 AVSS 0.724407f
C3208 a_n13990_8177.n14 AVSS 0.794542f
C3209 a_n13990_8177.n15 AVSS 0.542775f
C3210 a_n13990_8177.n16 AVSS 0.806162f
C3211 a_n13990_8177.n17 AVSS 0.806161f
C3212 a_n13990_8177.n18 AVSS 0.428083f
C3213 a_n13990_8177.n19 AVSS 0.724407f
C3214 a_n13990_8177.n20 AVSS 0.794542f
C3215 a_n13990_8177.n21 AVSS 0.946539f
C3216 a_n13990_8177.n22 AVSS 0.833972f
C3217 a_n13990_8177.n23 AVSS 0.724407f
C3218 a_n13990_8177.n24 AVSS 0.794542f
C3219 a_n13990_8177.n25 AVSS 0.542775f
C3220 a_n13990_8177.n26 AVSS 0.806162f
C3221 a_n13990_8177.n27 AVSS 0.806161f
C3222 a_n13990_8177.n28 AVSS 0.428083f
C3223 a_n13990_8177.n29 AVSS 0.724407f
C3224 a_n13990_8177.n30 AVSS 0.794542f
C3225 a_n13990_8177.n31 AVSS 0.946539f
C3226 a_n13990_8177.n32 AVSS 0.523557f
C3227 a_n13990_8177.n33 AVSS 0.842988f
C3228 a_n13990_8177.n34 AVSS 0.842981f
C3229 a_n13990_8177.n35 AVSS 0.820905f
C3230 a_n13990_8177.n36 AVSS 0.338474f
C3231 a_n13990_8177.n37 AVSS 0.842988f
C3232 a_n13990_8177.n38 AVSS 1.18777f
C3233 a_n13990_8177.n39 AVSS 1.05608f
C3234 a_n13990_8177.n40 AVSS 0.842988f
C3235 a_n13990_8177.n41 AVSS 0.842981f
C3236 a_n13990_8177.n42 AVSS 0.820905f
C3237 a_n13990_8177.n43 AVSS 0.338474f
C3238 a_n13990_8177.n44 AVSS 0.842988f
C3239 a_n13990_8177.n45 AVSS 1.18777f
C3240 a_n13990_8177.t177 AVSS 0.065937f
C3241 a_n13990_8177.t215 AVSS 0.173717f
C3242 a_n13990_8177.t187 AVSS 0.184972f
C3243 a_n13990_8177.n46 AVSS 0.591939f
C3244 a_n13990_8177.n47 AVSS 0.543506f
C3245 a_n13990_8177.t209 AVSS 0.173717f
C3246 a_n13990_8177.t199 AVSS 0.184972f
C3247 a_n13990_8177.n48 AVSS 0.702228f
C3248 a_n13990_8177.t128 AVSS 0.065937f
C3249 a_n13990_8177.t247 AVSS 0.065937f
C3250 a_n13990_8177.n49 AVSS 0.167319f
C3251 a_n13990_8177.t184 AVSS 0.065937f
C3252 a_n13990_8177.t174 AVSS 0.065937f
C3253 a_n13990_8177.n50 AVSS 0.180575f
C3254 a_n13990_8177.n51 AVSS 0.458299f
C3255 a_n13990_8177.n52 AVSS 0.381924f
C3256 a_n13990_8177.n53 AVSS 2.6775f
C3257 a_n13990_8177.n54 AVSS 2.73275f
C3258 a_n13990_8177.t196 AVSS 0.065937f
C3259 a_n13990_8177.t208 AVSS 0.065937f
C3260 a_n13990_8177.n55 AVSS 0.306918f
C3261 a_n13990_8177.t149 AVSS 0.298209f
C3262 a_n13990_8177.t255 AVSS 0.065937f
C3263 a_n13990_8177.t132 AVSS 0.065937f
C3264 a_n13990_8177.n56 AVSS 0.306918f
C3265 a_n13990_8177.t260 AVSS 0.5404f
C3266 a_n13990_8177.n57 AVSS 3.93851f
C3267 a_n13990_8177.t204 AVSS 0.065937f
C3268 a_n13990_8177.t258 AVSS 0.065937f
C3269 a_n13990_8177.n58 AVSS 0.633786f
C3270 a_n13990_8177.t213 AVSS 0.296468f
C3271 a_n13990_8177.n59 AVSS 1.70039f
C3272 a_n13990_8177.n60 AVSS 1.7652f
C3273 a_n13990_8177.t256 AVSS 0.065937f
C3274 a_n13990_8177.t137 AVSS 0.065937f
C3275 a_n13990_8177.n61 AVSS 0.304483f
C3276 a_n13990_8177.n62 AVSS 1.49371f
C3277 a_n13990_8177.t223 AVSS 0.296468f
C3278 a_n13990_8177.n63 AVSS 1.39244f
C3279 a_n13990_8177.t127 AVSS 0.173717f
C3280 a_n13990_8177.t138 AVSS 0.184972f
C3281 a_n13990_8177.n64 AVSS 0.702228f
C3282 a_n13990_8177.t233 AVSS 0.065937f
C3283 a_n13990_8177.t181 AVSS 0.065937f
C3284 a_n13990_8177.n65 AVSS 0.167319f
C3285 a_n13990_8177.t241 AVSS 0.065937f
C3286 a_n13990_8177.t191 AVSS 0.065937f
C3287 a_n13990_8177.n66 AVSS 0.180575f
C3288 a_n13990_8177.n67 AVSS 0.458299f
C3289 a_n13990_8177.n68 AVSS 0.381924f
C3290 a_n13990_8177.t253 AVSS 0.173717f
C3291 a_n13990_8177.t266 AVSS 0.184972f
C3292 a_n13990_8177.n69 AVSS 0.701534f
C3293 a_n13990_8177.t143 AVSS 0.065937f
C3294 a_n13990_8177.t262 AVSS 0.065937f
C3295 a_n13990_8177.n70 AVSS 0.167319f
C3296 a_n13990_8177.t152 AVSS 0.065937f
C3297 a_n13990_8177.t98 AVSS 0.065937f
C3298 a_n13990_8177.n71 AVSS 0.180575f
C3299 a_n13990_8177.n72 AVSS 0.458299f
C3300 a_n13990_8177.n73 AVSS 0.484178f
C3301 a_n13990_8177.t110 AVSS 0.173717f
C3302 a_n13990_8177.t116 AVSS 0.184972f
C3303 a_n13990_8177.n74 AVSS 0.583233f
C3304 a_n13990_8177.n75 AVSS 0.533851f
C3305 a_n13990_8177.t229 AVSS 0.173717f
C3306 a_n13990_8177.t234 AVSS 0.184972f
C3307 a_n13990_8177.n76 AVSS 0.585662f
C3308 a_n13990_8177.n77 AVSS 0.451282f
C3309 a_n13990_8177.n78 AVSS 0.181417f
C3310 a_n13990_8177.t243 AVSS 0.065937f
C3311 a_n13990_8177.t169 AVSS 0.065937f
C3312 a_n13990_8177.n79 AVSS 0.167319f
C3313 a_n13990_8177.t251 AVSS 0.065937f
C3314 a_n13990_8177.t178 AVSS 0.065937f
C3315 a_n13990_8177.n80 AVSS 0.180575f
C3316 a_n13990_8177.n81 AVSS 0.458299f
C3317 a_n13990_8177.n82 AVSS 0.25486f
C3318 a_n13990_8177.t190 AVSS 0.173717f
C3319 a_n13990_8177.t202 AVSS 0.184972f
C3320 a_n13990_8177.n83 AVSS 0.591939f
C3321 a_n13990_8177.n84 AVSS 0.543525f
C3322 a_n13990_8177.t134 AVSS 0.173717f
C3323 a_n13990_8177.t146 AVSS 0.184972f
C3324 a_n13990_8177.n85 AVSS 0.591939f
C3325 a_n13990_8177.n86 AVSS 0.543506f
C3326 a_n13990_8177.t155 AVSS 0.065937f
C3327 a_n13990_8177.t101 AVSS 0.065937f
C3328 a_n13990_8177.n87 AVSS 0.167319f
C3329 a_n13990_8177.t168 AVSS 0.065937f
C3330 a_n13990_8177.t113 AVSS 0.065937f
C3331 a_n13990_8177.n88 AVSS 0.180575f
C3332 a_n13990_8177.n89 AVSS 0.458299f
C3333 a_n13990_8177.n90 AVSS 0.357941f
C3334 a_n13990_8177.t119 AVSS 0.173717f
C3335 a_n13990_8177.t126 AVSS 0.184972f
C3336 a_n13990_8177.n91 AVSS 0.583233f
C3337 a_n13990_8177.n92 AVSS 0.533851f
C3338 a_n13990_8177.t185 AVSS 0.173717f
C3339 a_n13990_8177.t194 AVSS 0.184972f
C3340 a_n13990_8177.n93 AVSS 0.585662f
C3341 a_n13990_8177.n94 AVSS 0.451282f
C3342 a_n13990_8177.n95 AVSS 0.181417f
C3343 a_n13990_8177.n96 AVSS 4.29625f
C3344 a_n13990_8177.n97 AVSS 2.87631f
C3345 a_n13990_8177.t238 AVSS 0.065937f
C3346 a_n13990_8177.t107 AVSS 0.065937f
C3347 a_n13990_8177.n98 AVSS 0.306918f
C3348 a_n13990_8177.t163 AVSS 0.298209f
C3349 a_n13990_8177.t230 AVSS 0.065937f
C3350 a_n13990_8177.t225 AVSS 0.065937f
C3351 a_n13990_8177.n99 AVSS 0.306918f
C3352 a_n13990_8177.t109 AVSS 0.5404f
C3353 a_n13990_8177.n100 AVSS 1.25177f
C3354 a_n13990_8177.n101 AVSS 2.49893f
C3355 a_n13990_8177.t117 AVSS 0.296468f
C3356 a_n13990_8177.n102 AVSS 0.982185f
C3357 a_n13990_8177.t153 AVSS 0.065937f
C3358 a_n13990_8177.t216 AVSS 0.065937f
C3359 a_n13990_8177.n103 AVSS 0.304483f
C3360 a_n13990_8177.n104 AVSS 1.49371f
C3361 a_n13990_8177.t100 AVSS 0.065937f
C3362 a_n13990_8177.t156 AVSS 0.065937f
C3363 a_n13990_8177.n105 AVSS 0.633786f
C3364 a_n13990_8177.t108 AVSS 0.296468f
C3365 a_n13990_8177.n106 AVSS 1.70039f
C3366 a_n13990_8177.n107 AVSS 1.25245f
C3367 a_n13990_8177.n108 AVSS 2.42225f
C3368 a_n13990_8177.t259 AVSS 0.173717f
C3369 a_n13990_8177.t180 AVSS 0.184972f
C3370 a_n13990_8177.n109 AVSS 0.591939f
C3371 a_n13990_8177.n110 AVSS 0.543525f
C3372 a_n13990_8177.t140 AVSS 0.065937f
C3373 a_n13990_8177.t236 AVSS 0.065937f
C3374 a_n13990_8177.n111 AVSS 0.167319f
C3375 a_n13990_8177.t125 AVSS 0.065937f
C3376 a_n13990_8177.t268 AVSS 0.065937f
C3377 a_n13990_8177.n112 AVSS 0.180575f
C3378 a_n13990_8177.n113 AVSS 0.458299f
C3379 a_n13990_8177.n114 AVSS 0.25486f
C3380 a_n13990_8177.t151 AVSS 0.173717f
C3381 a_n13990_8177.t120 AVSS 0.184972f
C3382 a_n13990_8177.n115 AVSS 0.701534f
C3383 a_n13990_8177.t218 AVSS 0.065937f
C3384 a_n13990_8177.t159 AVSS 0.065937f
C3385 a_n13990_8177.n116 AVSS 0.167319f
C3386 a_n13990_8177.t160 AVSS 0.065937f
C3387 a_n13990_8177.t235 AVSS 0.065937f
C3388 a_n13990_8177.n117 AVSS 0.180575f
C3389 a_n13990_8177.n118 AVSS 0.458299f
C3390 a_n13990_8177.n119 AVSS 0.484178f
C3391 a_n13990_8177.t179 AVSS 0.173717f
C3392 a_n13990_8177.t147 AVSS 0.184972f
C3393 a_n13990_8177.n120 AVSS 0.583233f
C3394 a_n13990_8177.n121 AVSS 0.533851f
C3395 a_n13990_8177.t122 AVSS 0.173717f
C3396 a_n13990_8177.t220 AVSS 0.184972f
C3397 a_n13990_8177.n122 AVSS 0.585662f
C3398 a_n13990_8177.n123 AVSS 0.451282f
C3399 a_n13990_8177.n124 AVSS 0.181417f
C3400 a_n13990_8177.n125 AVSS 2.89625f
C3401 a_n13990_8177.n126 AVSS 2.52449f
C3402 a_n13990_8177.n127 AVSS 3.19912f
C3403 a_n13990_8177.t78 AVSS 0.260672f
C3404 a_n13990_8177.t19 AVSS 0.065937f
C3405 a_n13990_8177.t335 AVSS 0.065937f
C3406 a_n13990_8177.n128 AVSS 0.262999f
C3407 a_n13990_8177.t26 AVSS 0.260672f
C3408 a_n13990_8177.t291 AVSS 0.065937f
C3409 a_n13990_8177.t21 AVSS 0.065937f
C3410 a_n13990_8177.n129 AVSS 0.603414f
C3411 a_n13990_8177.t28 AVSS 0.260672f
C3412 a_n13990_8177.t29 AVSS 0.065937f
C3413 a_n13990_8177.t321 AVSS 0.065937f
C3414 a_n13990_8177.n130 AVSS 0.603414f
C3415 a_n13990_8177.n131 AVSS 1.7851f
C3416 a_n13990_8177.t35 AVSS 0.260672f
C3417 a_n13990_8177.t348 AVSS 0.065937f
C3418 a_n13990_8177.t342 AVSS 0.065937f
C3419 a_n13990_8177.n132 AVSS 0.262999f
C3420 a_n13990_8177.n133 AVSS 4.43096f
C3421 a_n13990_8177.t2 AVSS 0.065937f
C3422 a_n13990_8177.t45 AVSS 0.065937f
C3423 a_n13990_8177.n134 AVSS 0.197755f
C3424 a_n13990_8177.t4 AVSS 0.065937f
C3425 a_n13990_8177.t46 AVSS 0.065937f
C3426 a_n13990_8177.n135 AVSS 0.153269f
C3427 a_n13990_8177.n136 AVSS 0.455172f
C3428 a_n13990_8177.n137 AVSS 0.395084f
C3429 a_n13990_8177.t20 AVSS 0.065937f
C3430 a_n13990_8177.t17 AVSS 0.065937f
C3431 a_n13990_8177.n138 AVSS 0.197755f
C3432 a_n13990_8177.t12 AVSS 0.065937f
C3433 a_n13990_8177.t18 AVSS 0.065937f
C3434 a_n13990_8177.n139 AVSS 0.153269f
C3435 a_n13990_8177.n140 AVSS 0.455172f
C3436 a_n13990_8177.n141 AVSS 0.710232f
C3437 a_n13990_8177.t332 AVSS 0.065937f
C3438 a_n13990_8177.t10 AVSS 0.065937f
C3439 a_n13990_8177.n142 AVSS 0.197755f
C3440 a_n13990_8177.t334 AVSS 0.065937f
C3441 a_n13990_8177.t11 AVSS 0.065937f
C3442 a_n13990_8177.n143 AVSS 0.153269f
C3443 a_n13990_8177.n144 AVSS 0.455172f
C3444 a_n13990_8177.n145 AVSS 0.71025f
C3445 a_n13990_8177.t306 AVSS 0.065937f
C3446 a_n13990_8177.t343 AVSS 0.065937f
C3447 a_n13990_8177.n146 AVSS 0.197755f
C3448 a_n13990_8177.t317 AVSS 0.065937f
C3449 a_n13990_8177.t345 AVSS 0.065937f
C3450 a_n13990_8177.n147 AVSS 0.153269f
C3451 a_n13990_8177.n148 AVSS 0.455172f
C3452 a_n13990_8177.n149 AVSS 0.700453f
C3453 a_n13990_8177.t318 AVSS 0.065937f
C3454 a_n13990_8177.t347 AVSS 0.065937f
C3455 a_n13990_8177.n150 AVSS 0.197755f
C3456 a_n13990_8177.t319 AVSS 0.065937f
C3457 a_n13990_8177.t350 AVSS 0.065937f
C3458 a_n13990_8177.n151 AVSS 0.153269f
C3459 a_n13990_8177.n152 AVSS 0.63464f
C3460 a_n13990_8177.t81 AVSS 0.065937f
C3461 a_n13990_8177.t84 AVSS 0.065937f
C3462 a_n13990_8177.n153 AVSS 0.197755f
C3463 a_n13990_8177.t304 AVSS 0.065937f
C3464 a_n13990_8177.t85 AVSS 0.065937f
C3465 a_n13990_8177.n154 AVSS 0.153269f
C3466 a_n13990_8177.n155 AVSS 0.455172f
C3467 a_n13990_8177.n156 AVSS 0.917032f
C3468 a_n13990_8177.t8 AVSS 0.065937f
C3469 a_n13990_8177.t39 AVSS 0.065937f
C3470 a_n13990_8177.n157 AVSS 0.197755f
C3471 a_n13990_8177.t9 AVSS 0.065937f
C3472 a_n13990_8177.t41 AVSS 0.065937f
C3473 a_n13990_8177.n158 AVSS 0.153269f
C3474 a_n13990_8177.n159 AVSS 0.455172f
C3475 a_n13990_8177.n160 AVSS 0.710232f
C3476 a_n13990_8177.t23 AVSS 0.065937f
C3477 a_n13990_8177.t289 AVSS 0.065937f
C3478 a_n13990_8177.n161 AVSS 0.197755f
C3479 a_n13990_8177.t24 AVSS 0.065937f
C3480 a_n13990_8177.t290 AVSS 0.065937f
C3481 a_n13990_8177.n162 AVSS 0.153269f
C3482 a_n13990_8177.n163 AVSS 0.455172f
C3483 a_n13990_8177.n164 AVSS 0.188712f
C3484 a_n13990_8177.n165 AVSS 0.554552f
C3485 a_n13990_8177.n166 AVSS 3.89079f
C3486 a_n13990_8177.t22 AVSS 0.065937f
C3487 a_n13990_8177.t38 AVSS 0.065937f
C3488 a_n13990_8177.n167 AVSS 0.263575f
C3489 a_n13990_8177.n168 AVSS 0.962259f
C3490 a_n13990_8177.t80 AVSS 0.261154f
C3491 a_n13990_8177.n169 AVSS 1.24523f
C3492 a_n13990_8177.t37 AVSS 0.506358f
C3493 a_n13990_8177.t13 AVSS 0.065937f
C3494 a_n13990_8177.t16 AVSS 0.065937f
C3495 a_n13990_8177.n170 AVSS 0.263575f
C3496 a_n13990_8177.n171 AVSS 1.78417f
C3497 a_n13990_8177.n172 AVSS 1.25132f
C3498 a_n13990_8177.n173 AVSS 2.79169f
C3499 a_n13990_8177.n174 AVSS 2.50125f
C3500 a_n13990_8177.n175 AVSS 1.25252f
C3501 a_n13990_8177.n176 AVSS 2.77274f
C3502 a_n13990_8177.t31 AVSS 0.065937f
C3503 a_n13990_8177.t288 AVSS 0.065937f
C3504 a_n13990_8177.n177 AVSS 0.197755f
C3505 a_n13990_8177.t30 AVSS 0.065937f
C3506 a_n13990_8177.t351 AVSS 0.065937f
C3507 a_n13990_8177.n178 AVSS 0.153269f
C3508 a_n13990_8177.n179 AVSS 0.63464f
C3509 a_n13990_8177.t305 AVSS 0.065937f
C3510 a_n13990_8177.t79 AVSS 0.065937f
C3511 a_n13990_8177.n180 AVSS 0.197755f
C3512 a_n13990_8177.t303 AVSS 0.065937f
C3513 a_n13990_8177.t336 AVSS 0.065937f
C3514 a_n13990_8177.n181 AVSS 0.153269f
C3515 a_n13990_8177.n182 AVSS 0.455172f
C3516 a_n13990_8177.n183 AVSS 0.917032f
C3517 a_n13990_8177.t34 AVSS 0.065937f
C3518 a_n13990_8177.t7 AVSS 0.065937f
C3519 a_n13990_8177.n184 AVSS 0.197755f
C3520 a_n13990_8177.t33 AVSS 0.065937f
C3521 a_n13990_8177.t15 AVSS 0.065937f
C3522 a_n13990_8177.n185 AVSS 0.153269f
C3523 a_n13990_8177.n186 AVSS 0.455172f
C3524 a_n13990_8177.n187 AVSS 0.710232f
C3525 a_n13990_8177.t56 AVSS 0.065937f
C3526 a_n13990_8177.t349 AVSS 0.065937f
C3527 a_n13990_8177.n188 AVSS 0.197755f
C3528 a_n13990_8177.t55 AVSS 0.065937f
C3529 a_n13990_8177.t320 AVSS 0.065937f
C3530 a_n13990_8177.n189 AVSS 0.153269f
C3531 a_n13990_8177.n190 AVSS 0.455172f
C3532 a_n13990_8177.n191 AVSS 0.188712f
C3533 a_n13990_8177.n192 AVSS 0.554552f
C3534 a_n13990_8177.t3 AVSS 0.065937f
C3535 a_n13990_8177.t344 AVSS 0.065937f
C3536 a_n13990_8177.n193 AVSS 0.197755f
C3537 a_n13990_8177.t57 AVSS 0.065937f
C3538 a_n13990_8177.t86 AVSS 0.065937f
C3539 a_n13990_8177.n194 AVSS 0.153269f
C3540 a_n13990_8177.n195 AVSS 0.455172f
C3541 a_n13990_8177.n196 AVSS 0.700453f
C3542 a_n13990_8177.t27 AVSS 0.065937f
C3543 a_n13990_8177.t32 AVSS 0.065937f
C3544 a_n13990_8177.n197 AVSS 0.197755f
C3545 a_n13990_8177.t36 AVSS 0.065937f
C3546 a_n13990_8177.t40 AVSS 0.065937f
C3547 a_n13990_8177.n198 AVSS 0.153269f
C3548 a_n13990_8177.n199 AVSS 0.455172f
C3549 a_n13990_8177.n200 AVSS 0.71025f
C3550 a_n13990_8177.t6 AVSS 0.065937f
C3551 a_n13990_8177.t44 AVSS 0.065937f
C3552 a_n13990_8177.n201 AVSS 0.197755f
C3553 a_n13990_8177.t5 AVSS 0.065937f
C3554 a_n13990_8177.t43 AVSS 0.065937f
C3555 a_n13990_8177.n202 AVSS 0.153269f
C3556 a_n13990_8177.n203 AVSS 0.455172f
C3557 a_n13990_8177.n204 AVSS 0.710232f
C3558 a_n13990_8177.t83 AVSS 0.065937f
C3559 a_n13990_8177.t54 AVSS 0.065937f
C3560 a_n13990_8177.n205 AVSS 0.197755f
C3561 a_n13990_8177.t82 AVSS 0.065937f
C3562 a_n13990_8177.t346 AVSS 0.065937f
C3563 a_n13990_8177.n206 AVSS 0.153269f
C3564 a_n13990_8177.n207 AVSS 0.455172f
C3565 a_n13990_8177.n208 AVSS 0.395084f
C3566 a_n13990_8177.n209 AVSS 2.54508f
C3567 a_n13990_8177.n210 AVSS 3.86208f
C3568 a_n13990_8177.t14 AVSS 0.065937f
C3569 a_n13990_8177.t25 AVSS 0.065937f
C3570 a_n13990_8177.n211 AVSS 0.263575f
C3571 a_n13990_8177.n212 AVSS 0.962259f
C3572 a_n13990_8177.t53 AVSS 0.261154f
C3573 a_n13990_8177.n213 AVSS 1.24523f
C3574 a_n13990_8177.t292 AVSS 0.506358f
C3575 a_n13990_8177.t42 AVSS 0.065937f
C3576 a_n13990_8177.t333 AVSS 0.065937f
C3577 a_n13990_8177.n214 AVSS 0.263575f
C3578 a_n13990_8177.n215 AVSS 1.78417f
C3579 a_n13990_8177.n216 AVSS 1.25132f
C3580 a_n13990_8177.n217 AVSS 3.1335f
C3581 a_n13990_8177.n218 AVSS 2.00968f
C3582 a_n13990_8177.n219 AVSS 3.43055f
C3583 a_n13990_8177.n220 AVSS 3.1205f
C3584 a_n13990_8177.t182 AVSS 0.372643f
C3585 a_n13990_8177.t165 AVSS 0.065937f
C3586 a_n13990_8177.t157 AVSS 0.065937f
C3587 a_n13990_8177.n221 AVSS 0.284868f
C3588 a_n13990_8177.t269 AVSS 0.279265f
C3589 a_n13990_8177.t244 AVSS 0.278902f
C3590 a_n13990_8177.n222 AVSS 2.69004f
C3591 a_n13990_8177.t222 AVSS 0.369169f
C3592 a_n13990_8177.t145 AVSS 0.065937f
C3593 a_n13990_8177.t267 AVSS 0.065937f
C3594 a_n13990_8177.n223 AVSS 0.285448f
C3595 a_n13990_8177.n224 AVSS 0.939609f
C3596 a_n13990_8177.t270 AVSS 0.279833f
C3597 a_n13990_8177.n225 AVSS 0.79527f
C3598 a_n13990_8177.t212 AVSS 0.277438f
C3599 a_n13990_8177.n226 AVSS 0.720573f
C3600 a_n13990_8177.t170 AVSS 0.374369f
C3601 a_n13990_8177.t232 AVSS 0.065937f
C3602 a_n13990_8177.t176 AVSS 0.065937f
C3603 a_n13990_8177.n227 AVSS 0.285448f
C3604 a_n13990_8177.n228 AVSS 0.837957f
C3605 a_n13990_8177.t272 AVSS 0.374369f
C3606 a_n13990_8177.t161 AVSS 0.065937f
C3607 a_n13990_8177.t105 AVSS 0.065937f
C3608 a_n13990_8177.n229 AVSS 0.285448f
C3609 a_n13990_8177.n230 AVSS 0.837957f
C3610 a_n13990_8177.n231 AVSS 0.642415f
C3611 a_n13990_8177.t210 AVSS 0.162516f
C3612 a_n13990_8177.t217 AVSS 0.198291f
C3613 a_n13990_8177.n232 AVSS 1.06267f
C3614 a_n13990_8177.t239 AVSS 0.065937f
C3615 a_n13990_8177.t124 AVSS 0.065937f
C3616 a_n13990_8177.n233 AVSS 0.154318f
C3617 a_n13990_8177.t246 AVSS 0.065937f
C3618 a_n13990_8177.t130 AVSS 0.065937f
C3619 a_n13990_8177.n234 AVSS 0.196324f
C3620 a_n13990_8177.n235 AVSS 0.446846f
C3621 a_n13990_8177.n236 AVSS 0.976785f
C3622 a_n13990_8177.t144 AVSS 0.369169f
C3623 a_n13990_8177.t245 AVSS 0.065937f
C3624 a_n13990_8177.t198 AVSS 0.065937f
C3625 a_n13990_8177.n237 AVSS 0.285448f
C3626 a_n13990_8177.n238 AVSS 0.939609f
C3627 a_n13990_8177.t201 AVSS 0.279833f
C3628 a_n13990_8177.n239 AVSS 0.79527f
C3629 a_n13990_8177.t129 AVSS 0.277438f
C3630 a_n13990_8177.n240 AVSS 0.720573f
C3631 a_n13990_8177.t121 AVSS 0.277438f
C3632 a_n13990_8177.n241 AVSS 0.720573f
C3633 a_n13990_8177.t237 AVSS 0.279833f
C3634 a_n13990_8177.n242 AVSS 0.79527f
C3635 a_n13990_8177.t261 AVSS 0.065937f
C3636 a_n13990_8177.t186 AVSS 0.065937f
C3637 a_n13990_8177.n243 AVSS 0.285448f
C3638 a_n13990_8177.n244 AVSS 0.542568f
C3639 a_n13990_8177.t207 AVSS 0.277438f
C3640 a_n13990_8177.n245 AVSS 0.800289f
C3641 a_n13990_8177.t150 AVSS 0.279755f
C3642 a_n13990_8177.n246 AVSS 0.806849f
C3643 a_n13990_8177.t173 AVSS 0.065937f
C3644 a_n13990_8177.t115 AVSS 0.065937f
C3645 a_n13990_8177.n247 AVSS 0.285448f
C3646 a_n13990_8177.n248 AVSS 0.428365f
C3647 a_n13990_8177.n249 AVSS 0.642415f
C3648 a_n13990_8177.n250 AVSS 3.7876f
C3649 a_n13990_8177.n251 AVSS 1.2517f
C3650 a_n13990_8177.t193 AVSS 0.162516f
C3651 a_n13990_8177.t205 AVSS 0.198291f
C3652 a_n13990_8177.n252 AVSS 0.581115f
C3653 a_n13990_8177.n253 AVSS 1.18777f
C3654 a_n13990_8177.t188 AVSS 0.065937f
C3655 a_n13990_8177.t240 AVSS 0.065937f
C3656 a_n13990_8177.n254 AVSS 0.154318f
C3657 a_n13990_8177.t200 AVSS 0.065937f
C3658 a_n13990_8177.t249 AVSS 0.065937f
C3659 a_n13990_8177.n255 AVSS 0.196324f
C3660 a_n13990_8177.n256 AVSS 0.446846f
C3661 a_n13990_8177.n257 AVSS 0.776654f
C3662 a_n13990_8177.n258 AVSS 4.1989f
C3663 a_n13990_8177.t167 AVSS 0.372643f
C3664 a_n13990_8177.t271 AVSS 0.065937f
C3665 a_n13990_8177.t219 AVSS 0.065937f
C3666 a_n13990_8177.n259 AVSS 0.284868f
C3667 a_n13990_8177.t224 AVSS 0.279265f
C3668 a_n13990_8177.t154 AVSS 0.278902f
C3669 a_n13990_8177.n260 AVSS 0.183799f
C3670 a_n13990_8177.t195 AVSS 0.065937f
C3671 a_n13990_8177.t133 AVSS 0.065937f
C3672 a_n13990_8177.n261 AVSS 0.284868f
C3673 a_n13990_8177.t175 AVSS 0.279265f
C3674 a_n13990_8177.t226 AVSS 0.279265f
C3675 a_n13990_8177.t111 AVSS 0.065937f
C3676 a_n13990_8177.t211 AVSS 0.065937f
C3677 a_n13990_8177.n262 AVSS 0.284868f
C3678 a_n13990_8177.t263 AVSS 0.279265f
C3679 a_n13990_8177.t141 AVSS 0.278902f
C3680 a_n13990_8177.t183 AVSS 0.065937f
C3681 a_n13990_8177.t123 AVSS 0.065937f
C3682 a_n13990_8177.n263 AVSS 0.284868f
C3683 a_n13990_8177.t118 AVSS 0.373142f
C3684 a_n13990_8177.n264 AVSS 0.183799f
C3685 a_n13990_8177.n265 AVSS 2.69004f
C3686 a_n13990_8177.n266 AVSS 2.41819f
C3687 a_n13990_8177.n267 AVSS 0.183807f
C3688 a_n13990_8177.t197 AVSS 0.277438f
C3689 a_n13990_8177.n268 AVSS 0.720573f
C3690 a_n13990_8177.t135 AVSS 0.279833f
C3691 a_n13990_8177.n269 AVSS 0.79527f
C3692 a_n13990_8177.t158 AVSS 0.065937f
C3693 a_n13990_8177.t252 AVSS 0.065937f
C3694 a_n13990_8177.n270 AVSS 0.285448f
C3695 a_n13990_8177.n271 AVSS 0.542568f
C3696 a_n13990_8177.t102 AVSS 0.277438f
C3697 a_n13990_8177.n272 AVSS 0.800289f
C3698 a_n13990_8177.t228 AVSS 0.279755f
C3699 a_n13990_8177.n273 AVSS 0.806849f
C3700 a_n13990_8177.t242 AVSS 0.065937f
C3701 a_n13990_8177.t189 AVSS 0.065937f
C3702 a_n13990_8177.n274 AVSS 0.285448f
C3703 a_n13990_8177.n275 AVSS 0.428365f
C3704 a_n13990_8177.n276 AVSS 0.183807f
C3705 a_n13990_8177.n277 AVSS 2.41819f
C3706 a_n13990_8177.t104 AVSS 0.162516f
C3707 a_n13990_8177.t214 AVSS 0.198291f
C3708 a_n13990_8177.n278 AVSS 1.06267f
C3709 a_n13990_8177.t136 AVSS 0.065937f
C3710 a_n13990_8177.t203 AVSS 0.065937f
C3711 a_n13990_8177.n279 AVSS 0.154318f
C3712 a_n13990_8177.t221 AVSS 0.065937f
C3713 a_n13990_8177.t166 AVSS 0.065937f
C3714 a_n13990_8177.n280 AVSS 0.196324f
C3715 a_n13990_8177.n281 AVSS 0.446846f
C3716 a_n13990_8177.n282 AVSS 0.976785f
C3717 a_n13990_8177.t257 AVSS 0.065937f
C3718 a_n13990_8177.t139 AVSS 0.065937f
C3719 a_n13990_8177.n283 AVSS 0.154318f
C3720 a_n13990_8177.t148 AVSS 0.065937f
C3721 a_n13990_8177.t103 AVSS 0.065937f
C3722 a_n13990_8177.n284 AVSS 0.196324f
C3723 a_n13990_8177.n285 AVSS 0.446846f
C3724 a_n13990_8177.n286 AVSS 0.776654f
C3725 a_n13990_8177.t265 AVSS 0.162516f
C3726 a_n13990_8177.t99 AVSS 0.198291f
C3727 a_n13990_8177.n287 AVSS 0.581115f
C3728 a_n13990_8177.n288 AVSS 1.18777f
C3729 a_n13990_8177.n289 AVSS 1.2517f
C3730 a_n13990_8177.n290 AVSS 2.70921f
C3731 a_n13990_8177.n291 AVSS 2.6883f
C3732 a_n13990_8177.t66 AVSS 0.065937f
C3733 a_n13990_8177.t89 AVSS 0.065937f
C3734 a_n13990_8177.n292 AVSS 0.181906f
C3735 a_n13990_8177.t64 AVSS 0.065937f
C3736 a_n13990_8177.t87 AVSS 0.065937f
C3737 a_n13990_8177.n293 AVSS 0.166113f
C3738 a_n13990_8177.n294 AVSS 1.02196f
C3739 a_n13990_8177.t72 AVSS 0.186098f
C3740 a_n13990_8177.t70 AVSS 0.172688f
C3741 a_n13990_8177.n295 AVSS 0.591849f
C3742 a_n13990_8177.n296 AVSS 1.17271f
C3743 a_n13990_8177.n297 AVSS 4.22418f
C3744 a_n13990_8177.t60 AVSS 0.065937f
C3745 a_n13990_8177.t337 AVSS 0.065937f
C3746 a_n13990_8177.n298 AVSS 0.362252f
C3747 a_n13990_8177.t91 AVSS 0.065937f
C3748 a_n13990_8177.t90 AVSS 0.065937f
C3749 a_n13990_8177.n299 AVSS 0.241904f
C3750 a_n13990_8177.n300 AVSS 1.18973f
C3751 a_n13990_8177.t0 AVSS 0.065937f
C3752 a_n13990_8177.t314 AVSS 0.065937f
C3753 a_n13990_8177.n301 AVSS 0.241904f
C3754 a_n13990_8177.n302 AVSS 0.843783f
C3755 a_n13990_8177.t327 AVSS 0.065937f
C3756 a_n13990_8177.t69 AVSS 0.065937f
C3757 a_n13990_8177.n303 AVSS 0.241904f
C3758 a_n13990_8177.n304 AVSS 0.338896f
C3759 a_n13990_8177.t313 AVSS 0.065937f
C3760 a_n13990_8177.t274 AVSS 0.065937f
C3761 a_n13990_8177.n305 AVSS 0.361324f
C3762 a_n13990_8177.t296 AVSS 0.065937f
C3763 a_n13990_8177.t295 AVSS 0.065937f
C3764 a_n13990_8177.n306 AVSS 0.241201f
C3765 a_n13990_8177.t49 AVSS 0.065937f
C3766 a_n13990_8177.t88 AVSS 0.065937f
C3767 a_n13990_8177.n307 AVSS 0.241201f
C3768 a_n13990_8177.t62 AVSS 0.065937f
C3769 a_n13990_8177.t324 AVSS 0.065937f
C3770 a_n13990_8177.n308 AVSS 0.241201f
C3771 a_n13990_8177.t294 AVSS 0.065937f
C3772 a_n13990_8177.t328 AVSS 0.065937f
C3773 a_n13990_8177.n309 AVSS 0.241201f
C3774 a_n13990_8177.t74 AVSS 0.065937f
C3775 a_n13990_8177.t310 AVSS 0.065937f
C3776 a_n13990_8177.n310 AVSS 0.241201f
C3777 a_n13990_8177.t71 AVSS 0.065937f
C3778 a_n13990_8177.t67 AVSS 0.065937f
C3779 a_n13990_8177.n311 AVSS 0.241201f
C3780 a_n13990_8177.t47 AVSS 0.065937f
C3781 a_n13990_8177.t280 AVSS 0.065937f
C3782 a_n13990_8177.n312 AVSS 0.241201f
C3783 a_n13990_8177.n313 AVSS 1.13487f
C3784 a_n13990_8177.t340 AVSS 0.065937f
C3785 a_n13990_8177.t278 AVSS 0.065937f
C3786 a_n13990_8177.n314 AVSS 0.181906f
C3787 a_n13990_8177.t293 AVSS 0.065937f
C3788 a_n13990_8177.t309 AVSS 0.065937f
C3789 a_n13990_8177.n315 AVSS 0.166113f
C3790 a_n13990_8177.n316 AVSS 1.02196f
C3791 a_n13990_8177.t52 AVSS 0.186098f
C3792 a_n13990_8177.t68 AVSS 0.172688f
C3793 a_n13990_8177.n317 AVSS 0.591849f
C3794 a_n13990_8177.n318 AVSS 1.17271f
C3795 a_n13990_8177.t277 AVSS 0.186098f
C3796 a_n13990_8177.t307 AVSS 0.172688f
C3797 a_n13990_8177.n319 AVSS 0.591849f
C3798 a_n13990_8177.n320 AVSS 0.708323f
C3799 a_n13990_8177.t297 AVSS 0.065937f
C3800 a_n13990_8177.t285 AVSS 0.065937f
C3801 a_n13990_8177.n321 AVSS 0.181906f
C3802 a_n13990_8177.t283 AVSS 0.065937f
C3803 a_n13990_8177.t287 AVSS 0.065937f
C3804 a_n13990_8177.n322 AVSS 0.166113f
C3805 a_n13990_8177.n323 AVSS 0.458182f
C3806 a_n13990_8177.n324 AVSS 1.08733f
C3807 a_n13990_8177.n325 AVSS 1.25142f
C3808 a_n13990_8177.n326 AVSS 3.83833f
C3809 a_n13990_8177.n327 AVSS 2.79169f
C3810 a_n13990_8177.n328 AVSS 0.549878f
C3811 a_n13990_8177.t77 AVSS 0.065937f
C3812 a_n13990_8177.t96 AVSS 0.065937f
C3813 a_n13990_8177.n329 AVSS 0.241904f
C3814 a_n13990_8177.n330 AVSS 0.822008f
C3815 a_n13990_8177.t322 AVSS 0.065937f
C3816 a_n13990_8177.t338 AVSS 0.065937f
C3817 a_n13990_8177.n331 AVSS 0.241904f
C3818 a_n13990_8177.n332 AVSS 0.843765f
C3819 a_n13990_8177.t281 AVSS 0.065937f
C3820 a_n13990_8177.t50 AVSS 0.065937f
C3821 a_n13990_8177.n333 AVSS 0.241904f
C3822 a_n13990_8177.n334 AVSS 0.843783f
C3823 a_n13990_8177.t276 AVSS 0.065937f
C3824 a_n13990_8177.t308 AVSS 0.065937f
C3825 a_n13990_8177.n335 AVSS 0.241904f
C3826 a_n13990_8177.n336 AVSS 0.518837f
C3827 a_n13990_8177.n337 AVSS 2.81995f
C3828 a_n13990_8177.t95 AVSS 0.065937f
C3829 a_n13990_8177.t76 AVSS 0.065937f
C3830 a_n13990_8177.n338 AVSS 0.361324f
C3831 a_n13990_8177.t275 AVSS 0.065937f
C3832 a_n13990_8177.t315 AVSS 0.065937f
C3833 a_n13990_8177.n339 AVSS 0.241201f
C3834 a_n13990_8177.t61 AVSS 0.065937f
C3835 a_n13990_8177.t75 AVSS 0.065937f
C3836 a_n13990_8177.n340 AVSS 0.241201f
C3837 a_n13990_8177.t63 AVSS 0.065937f
C3838 a_n13990_8177.t97 AVSS 0.065937f
C3839 a_n13990_8177.n341 AVSS 0.241201f
C3840 a_n13990_8177.n342 AVSS 0.549825f
C3841 a_n13990_8177.t341 AVSS 0.065937f
C3842 a_n13990_8177.t316 AVSS 0.065937f
C3843 a_n13990_8177.n343 AVSS 0.241201f
C3844 a_n13990_8177.t329 AVSS 0.065937f
C3845 a_n13990_8177.t284 AVSS 0.065937f
C3846 a_n13990_8177.n344 AVSS 0.241201f
C3847 a_n13990_8177.t73 AVSS 0.065937f
C3848 a_n13990_8177.t331 AVSS 0.065937f
C3849 a_n13990_8177.n345 AVSS 0.241201f
C3850 a_n13990_8177.t94 AVSS 0.065937f
C3851 a_n13990_8177.t59 AVSS 0.065937f
C3852 a_n13990_8177.n346 AVSS 0.241201f
C3853 a_n13990_8177.n347 AVSS 2.71764f
C3854 a_n13990_8177.n348 AVSS 2.64144f
C3855 a_n13990_8177.t300 AVSS 0.186098f
C3856 a_n13990_8177.t299 AVSS 0.172688f
C3857 a_n13990_8177.n349 AVSS 0.591849f
C3858 a_n13990_8177.n350 AVSS 0.708322f
C3859 a_n13990_8177.t302 AVSS 0.065937f
C3860 a_n13990_8177.t92 AVSS 0.065937f
C3861 a_n13990_8177.n351 AVSS 0.181906f
C3862 a_n13990_8177.t301 AVSS 0.065937f
C3863 a_n13990_8177.t1 AVSS 0.065937f
C3864 a_n13990_8177.n352 AVSS 0.166113f
C3865 a_n13990_8177.n353 AVSS 0.458182f
C3866 a_n13990_8177.n354 AVSS 1.08733f
C3867 a_n13990_8177.n355 AVSS 1.25142f
C3868 a_n13990_8177.n356 AVSS 2.33745f
C3869 a_n13990_8177.t65 AVSS 0.065937f
C3870 a_n13990_8177.t325 AVSS 0.065937f
C3871 a_n13990_8177.n357 AVSS 0.362252f
C3872 a_n13990_8177.t48 AVSS 0.065937f
C3873 a_n13990_8177.t330 AVSS 0.065937f
C3874 a_n13990_8177.n358 AVSS 0.241904f
C3875 a_n13990_8177.n359 AVSS 1.18973f
C3876 a_n13990_8177.t298 AVSS 0.065937f
C3877 a_n13990_8177.t311 AVSS 0.065937f
C3878 a_n13990_8177.n360 AVSS 0.241904f
C3879 a_n13990_8177.n361 AVSS 0.843783f
C3880 a_n13990_8177.t312 AVSS 0.065937f
C3881 a_n13990_8177.t323 AVSS 0.065937f
C3882 a_n13990_8177.n362 AVSS 0.241904f
C3883 a_n13990_8177.n363 AVSS 0.338896f
C3884 a_n13990_8177.t339 AVSS 0.065937f
C3885 a_n13990_8177.t282 AVSS 0.065937f
C3886 a_n13990_8177.n364 AVSS 0.241904f
C3887 a_n13990_8177.n365 AVSS 0.518837f
C3888 a_n13990_8177.t58 AVSS 0.065937f
C3889 a_n13990_8177.t51 AVSS 0.065937f
C3890 a_n13990_8177.n366 AVSS 0.241904f
C3891 a_n13990_8177.n367 AVSS 0.843783f
C3892 a_n13990_8177.t93 AVSS 0.065937f
C3893 a_n13990_8177.t286 AVSS 0.065937f
C3894 a_n13990_8177.n368 AVSS 0.241904f
C3895 a_n13990_8177.n369 AVSS 0.843765f
C3896 a_n13990_8177.t326 AVSS 0.065937f
C3897 a_n13990_8177.t279 AVSS 0.065937f
C3898 a_n13990_8177.n370 AVSS 0.241904f
C3899 a_n13990_8177.n371 AVSS 0.822008f
C3900 a_n13990_8177.n372 AVSS 0.549878f
C3901 a_n13990_8177.n373 AVSS 3.07641f
C3902 a_n13990_8177.n374 AVSS 2.08409f
C3903 a_n13990_8177.n375 AVSS 2.09974f
C3904 a_n13990_8177.n376 AVSS 3.0578f
C3905 a_n13990_8177.n377 AVSS 0.183799f
C3906 a_n13990_8177.t254 AVSS 0.065937f
C3907 a_n13990_8177.t162 AVSS 0.065937f
C3908 a_n13990_8177.n378 AVSS 0.284868f
C3909 a_n13990_8177.t171 AVSS 0.279265f
C3910 a_n13990_8177.t164 AVSS 0.279265f
C3911 a_n13990_8177.t114 AVSS 0.065937f
C3912 a_n13990_8177.t248 AVSS 0.065937f
C3913 a_n13990_8177.n379 AVSS 0.284868f
C3914 a_n13990_8177.t206 AVSS 0.279265f
C3915 a_n13990_8177.t131 AVSS 0.278902f
C3916 a_n13990_8177.t142 AVSS 0.065937f
C3917 a_n13990_8177.t227 AVSS 0.065937f
C3918 a_n13990_8177.n380 AVSS 0.284868f
C3919 a_n13990_8177.t106 AVSS 0.373142f
C3920 a_n13990_8177.n381 AVSS 0.183799f
C3921 a_n13990_8177.n382 AVSS 3.04283f
C3922 a_n13990_8177.n383 AVSS 2.84217f
C3923 a_n13990_8177.n384 AVSS 2.10814f
C3924 a_n13990_8177.n385 AVSS 2.84853f
C3925 a_n13990_8177.n386 AVSS 1.25177f
C3926 a_n13990_8177.n387 AVSS 3.2993f
C3927 a_n13990_8177.n388 AVSS 2.89625f
C3928 a_n13990_8177.n389 AVSS 0.181417f
C3929 a_n13990_8177.t250 AVSS 0.173717f
C3930 a_n13990_8177.t112 AVSS 0.184972f
C3931 a_n13990_8177.n390 AVSS 0.585662f
C3932 a_n13990_8177.n391 AVSS 0.451282f
C3933 a_n13990_8177.t192 AVSS 0.173717f
C3934 a_n13990_8177.t264 AVSS 0.184972f
C3935 a_n13990_8177.n392 AVSS 0.583233f
C3936 a_n13990_8177.n393 AVSS 0.533851f
C3937 a_n13990_8177.n394 AVSS 0.357941f
C3938 a_n13990_8177.t231 AVSS 0.065937f
C3939 a_n13990_8177.t172 AVSS 0.065937f
C3940 a_n13990_8177.n395 AVSS 0.167319f
C3941 a_n13990_8177.n396 AVSS 0.458299f
C3942 a_n13990_8177.n397 AVSS 0.180575f
C3943 a_n13990_8177.t273 AVSS 0.065937f
C3944 a_n11737_n15980.n0 AVSS 0.20217f
C3945 a_n11737_n15980.n1 AVSS 0.079131f
C3946 a_n11737_n15980.n2 AVSS 0.09668f
C3947 a_n11737_n15980.n3 AVSS 0.634055f
C3948 a_n11737_n15980.n4 AVSS 0.138006f
C3949 a_n11737_n15980.n5 AVSS 0.19395f
C3950 a_n11737_n15980.n6 AVSS 0.105198f
C3951 a_n11737_n15980.n7 AVSS 0.601785f
C3952 a_n11737_n15980.n8 AVSS 0.114218f
C3953 a_n11737_n15980.n9 AVSS 0.109304f
C3954 a_n11737_n15980.n10 AVSS 0.096682f
C3955 a_n11737_n15980.n11 AVSS 0.630679f
C3956 a_n11737_n15980.n12 AVSS 0.137093f
C3957 a_n11737_n15980.n13 AVSS 0.636534f
C3958 a_n11737_n15980.n14 AVSS 0.138019f
C3959 a_n11737_n15980.n15 AVSS 0.19088f
C3960 a_n11737_n15980.n16 AVSS 0.073662f
C3961 a_n11737_n15980.n17 AVSS 0.620893f
C3962 a_n11737_n15980.n18 AVSS 0.115211f
C3963 a_n11737_n15980.n19 AVSS 0.109353f
C3964 a_n11737_n15980.n20 AVSS 0.091177f
C3965 a_n11737_n15980.n21 AVSS 0.60394f
C3966 a_n11737_n15980.n22 AVSS 0.137085f
C3967 a_n11737_n15980.n23 AVSS 0.142063f
C3968 a_n11737_n15980.n24 AVSS 0.142376f
C3969 a_n11737_n15980.n25 AVSS 0.572195f
C3970 a_n11737_n15980.n26 AVSS 0.223163f
C3971 a_n11737_n15980.n27 AVSS 0.085766f
C3972 a_n11737_n15980.n28 AVSS 0.125036f
C3973 a_n11737_n15980.n29 AVSS 0.028544f
C3974 a_n11737_n15980.n30 AVSS 0.128752f
C3975 a_n11737_n15980.n31 AVSS 0.079498f
C3976 a_n11737_n15980.n32 AVSS 0.139663f
C3977 a_n11737_n15980.n33 AVSS 0.059501f
C3978 a_n11737_n15980.n34 AVSS 0.367432f
C3979 a_n11737_n15980.n35 AVSS 0.219253f
C3980 a_n11737_n15980.n36 AVSS 0.121627f
C3981 a_n11737_n15980.n37 AVSS 0.08337f
C3982 a_n11737_n15980.n38 AVSS 0.103678f
C3983 a_n11737_n15980.n39 AVSS 0.071374f
C3984 a_n11737_n15980.n40 AVSS 0.117473f
C3985 a_n11737_n15980.n41 AVSS 0.083871f
C3986 a_n11737_n15980.t11 AVSS 0.139831f
C3987 a_n11737_n15980.t22 AVSS 0.138588f
C3988 a_n11737_n15980.n42 AVSS 0.225221f
C3989 a_n11737_n15980.n43 AVSS 0.028243f
C3990 a_n11737_n15980.t5 AVSS 0.069996f
C3991 a_n11737_n15980.t7 AVSS 0.070436f
C3992 a_n11737_n15980.t13 AVSS 0.14362f
C3993 a_n11737_n15980.t18 AVSS 0.027525f
C3994 a_n11737_n15980.t6 AVSS 0.027525f
C3995 a_n11737_n15980.n44 AVSS 0.106569f
C3996 a_n11737_n15980.n45 AVSS 0.366596f
C3997 a_n11737_n15980.t15 AVSS 0.106099f
C3998 a_n11737_n15980.n46 AVSS 0.223009f
C3999 a_n11737_n15980.t3 AVSS 0.027525f
C4000 a_n11737_n15980.t2 AVSS 0.027525f
C4001 a_n11737_n15980.n47 AVSS 0.107073f
C4002 a_n11737_n15980.n48 AVSS 0.189205f
C4003 a_n11737_n15980.n49 AVSS 0.011282f
C4004 a_n11737_n15980.n50 AVSS 0.117789f
C4005 a_n11737_n15980.n51 AVSS 0.077478f
C4006 a_n11737_n15980.t10 AVSS 0.027525f
C4007 a_n11737_n15980.t9 AVSS 0.027525f
C4008 a_n11737_n15980.n52 AVSS 0.066904f
C4009 a_n11737_n15980.n53 AVSS 0.102145f
C4010 a_n11737_n15980.n54 AVSS 0.066599f
C4011 a_n11737_n15980.n55 AVSS 0.719637f
C4012 a_n11737_n15980.t44 AVSS 0.170059f
C4013 a_n11737_n15980.t27 AVSS 0.170823f
C4014 a_n11737_n15980.n56 AVSS 0.293789f
C4015 a_n11737_n15980.t48 AVSS 0.170054f
C4016 a_n11737_n15980.t36 AVSS 0.170854f
C4017 a_n11737_n15980.n57 AVSS 0.283517f
C4018 a_n11737_n15980.n58 AVSS 0.460971f
C4019 a_n11737_n15980.t63 AVSS 0.170054f
C4020 a_n11737_n15980.t1 AVSS 0.039658f
C4021 a_n11737_n15980.t0 AVSS 0.148789f
C4022 a_n11737_n15980.n59 AVSS 0.166098f
C4023 a_n11737_n15980.n60 AVSS 0.200097f
C4024 a_n11737_n15980.n61 AVSS 0.35548f
C4025 a_n11737_n15980.t52 AVSS 0.228597f
C4026 a_n11737_n15980.n62 AVSS 0.190527f
C4027 a_n11737_n15980.n63 AVSS 0.136818f
C4028 a_n11737_n15980.t34 AVSS 0.228597f
C4029 a_n11737_n15980.n64 AVSS 0.138255f
C4030 a_n11737_n15980.t64 AVSS 0.228597f
C4031 a_n11737_n15980.t35 AVSS 0.228597f
C4032 a_n11737_n15980.n65 AVSS 0.081746f
C4033 a_n11737_n15980.n66 AVSS 0.066252f
C4034 a_n11737_n15980.t40 AVSS 0.228597f
C4035 a_n11737_n15980.t53 AVSS 0.228597f
C4036 a_n11737_n15980.t41 AVSS 0.228597f
C4037 a_n11737_n15980.t28 AVSS 0.228597f
C4038 a_n11737_n15980.t42 AVSS 0.228597f
C4039 a_n11737_n15980.n67 AVSS 0.028542f
C4040 a_n11737_n15980.n68 AVSS 0.076654f
C4041 a_n11737_n15980.n69 AVSS 0.146583f
C4042 a_n11737_n15980.t25 AVSS 0.228597f
C4043 a_n11737_n15980.n70 AVSS 0.184236f
C4044 a_n11737_n15980.n71 AVSS 0.138285f
C4045 a_n11737_n15980.t37 AVSS 0.228597f
C4046 a_n11737_n15980.t49 AVSS 0.228597f
C4047 a_n11737_n15980.n72 AVSS 0.138297f
C4048 a_n11737_n15980.t50 AVSS 0.228597f
C4049 a_n11737_n15980.n73 AVSS 0.081788f
C4050 a_n11737_n15980.n74 AVSS 0.066232f
C4051 a_n11737_n15980.t58 AVSS 0.228597f
C4052 a_n11737_n15980.t26 AVSS 0.228597f
C4053 a_n11737_n15980.t45 AVSS 0.228597f
C4054 a_n11737_n15980.n75 AVSS 0.142075f
C4055 a_n11737_n15980.t55 AVSS 0.228597f
C4056 a_n11737_n15980.n76 AVSS 0.126499f
C4057 a_n11737_n15980.n77 AVSS 0.080408f
C4058 a_n11737_n15980.t54 AVSS 0.228597f
C4059 a_n11737_n15980.n78 AVSS 2.42396f
C4060 a_n11737_n15980.n79 AVSS 0.135659f
C4061 a_n11737_n15980.n80 AVSS 0.023596f
C4062 a_n11737_n15980.n81 AVSS 0.122783f
C4063 a_n11737_n15980.t56 AVSS 0.232075f
C4064 a_n11737_n15980.n82 AVSS 0.177208f
C4065 a_n11737_n15980.t43 AVSS 0.228597f
C4066 a_n11737_n15980.n83 AVSS 0.11235f
C4067 a_n11737_n15980.n84 AVSS 0.009526f
C4068 a_n11737_n15980.n85 AVSS 0.023596f
C4069 a_n11737_n15980.n86 AVSS 0.024838f
C4070 a_n11737_n15980.n87 AVSS 0.024838f
C4071 a_n11737_n15980.n88 AVSS 0.016253f
C4072 a_n11737_n15980.n89 AVSS 0.009463f
C4073 a_n11737_n15980.t57 AVSS 0.228597f
C4074 a_n11737_n15980.n90 AVSS 0.088453f
C4075 a_n11737_n15980.n91 AVSS 0.07798f
C4076 a_n11737_n15980.t31 AVSS 0.228597f
C4077 a_n11737_n15980.n92 AVSS 0.186542f
C4078 a_n11737_n15980.t60 AVSS 0.228597f
C4079 a_n11737_n15980.n93 AVSS 0.150463f
C4080 a_n11737_n15980.t32 AVSS 0.228597f
C4081 a_n11737_n15980.n94 AVSS 0.185296f
C4082 a_n11737_n15980.n95 AVSS 0.026771f
C4083 a_n11737_n15980.t62 AVSS 0.233855f
C4084 a_n11737_n15980.t51 AVSS 0.228597f
C4085 a_n11737_n15980.n96 AVSS 0.117059f
C4086 a_n11737_n15980.n97 AVSS 0.195606f
C4087 a_n11737_n15980.n98 AVSS 0.147771f
C4088 a_n11737_n15980.t61 AVSS 0.228597f
C4089 a_n11737_n15980.n99 AVSS 0.624753f
C4090 a_n11737_n15980.n100 AVSS 0.134349f
C4091 a_n11737_n15980.n101 AVSS 0.016253f
C4092 a_n11737_n15980.n102 AVSS 0.027643f
C4093 a_n11737_n15980.t29 AVSS 0.233737f
C4094 a_n11737_n15980.n103 AVSS 0.191045f
C4095 a_n11737_n15980.t59 AVSS 0.228597f
C4096 a_n11737_n15980.n104 AVSS 0.116872f
C4097 a_n11737_n15980.n105 AVSS 0.026647f
C4098 a_n11737_n15980.n106 AVSS 0.134119f
C4099 a_n11737_n15980.n107 AVSS 0.029098f
C4100 a_n11737_n15980.n108 AVSS 0.016253f
C4101 a_n11737_n15980.n109 AVSS 0.008218f
C4102 a_n11737_n15980.t30 AVSS 0.228597f
C4103 a_n11737_n15980.n110 AVSS 0.088453f
C4104 a_n11737_n15980.n111 AVSS 0.077901f
C4105 a_n11737_n15980.t46 AVSS 0.228597f
C4106 a_n11737_n15980.n112 AVSS 0.186293f
C4107 a_n11737_n15980.t33 AVSS 0.228597f
C4108 a_n11737_n15980.n113 AVSS 0.15138f
C4109 a_n11737_n15980.t47 AVSS 0.228597f
C4110 a_n11737_n15980.n114 AVSS 0.184354f
C4111 a_n11737_n15980.n115 AVSS 0.027643f
C4112 a_n11737_n15980.t39 AVSS 0.232075f
C4113 a_n11737_n15980.n116 AVSS 0.18242f
C4114 a_n11737_n15980.t24 AVSS 0.228597f
C4115 a_n11737_n15980.n117 AVSS 0.11136f
C4116 a_n11737_n15980.n118 AVSS 0.008716f
C4117 a_n11737_n15980.n119 AVSS 0.1266f
C4118 a_n11737_n15980.n120 AVSS 0.029098f
C4119 a_n11737_n15980.n121 AVSS 0.029098f
C4120 a_n11737_n15980.n122 AVSS 0.026149f
C4121 a_n11737_n15980.t38 AVSS 0.228597f
C4122 a_n11737_n15980.n123 AVSS 0.088453f
C4123 a_n11737_n15980.n124 AVSS 0.009214f
C4124 a_n11737_n15980.n125 AVSS 0.076354f
C4125 a_n11737_n15980.n126 AVSS 0.049938f
C4126 a_n11737_n15980.n127 AVSS 0.168034f
C4127 a_n11737_n15980.n128 AVSS 2.24469f
C4128 a_n11737_n15980.n129 AVSS 4.68353f
C4129 a_n11737_n15980.n130 AVSS 4.47196f
C4130 a_n11737_n15980.n131 AVSS 2.60408f
C4131 a_n11737_n15980.n132 AVSS 0.01577f
C4132 a_n11737_n15980.n133 AVSS 0.226586f
C4133 a_n11737_n15980.t17 AVSS 0.027525f
C4134 a_n11737_n15980.t16 AVSS 0.027525f
C4135 a_n11737_n15980.n134 AVSS 0.067484f
C4136 a_n11737_n15980.t12 AVSS 0.1069f
C4137 a_n11737_n15980.t4 AVSS 0.027525f
C4138 a_n11737_n15980.t21 AVSS 0.027525f
C4139 a_n11737_n15980.n135 AVSS 0.106456f
C4140 a_n11737_n15980.n136 AVSS 0.187719f
C4141 a_n11737_n15980.n137 AVSS 0.081766f
C4142 a_n11737_n15980.t19 AVSS 0.070025f
C4143 a_n11737_n15980.n138 AVSS 0.1181f
C4144 a_n11737_n15980.n139 AVSS 0.011282f
C4145 a_n11737_n15980.n140 AVSS 0.02713f
C4146 a_n11737_n15980.t8 AVSS 0.027525f
C4147 a_n11737_n15980.t14 AVSS 0.027525f
C4148 a_n11737_n15980.n141 AVSS 0.107515f
C4149 a_n11737_n15980.t20 AVSS 0.144635f
C4150 a_n11737_n15980.t23 AVSS 0.070407f
C4151 IREF.t15 AVSS 0.046573f
C4152 IREF.t27 AVSS 0.046573f
C4153 IREF.n0 AVSS 0.111955f
C4154 IREF.n1 AVSS 0.061105f
C4155 IREF.n2 AVSS 0.0275f
C4156 IREF.n3 AVSS 0.0275f
C4157 IREF.n4 AVSS 0.0275f
C4158 IREF.t19 AVSS 0.23889f
C4159 IREF.n5 AVSS 0.386586f
C4160 IREF.t37 AVSS 0.046573f
C4161 IREF.t31 AVSS 0.046573f
C4162 IREF.n6 AVSS 0.115949f
C4163 IREF.n7 AVSS 0.118885f
C4164 IREF.n8 AVSS 0.061105f
C4165 IREF.n9 AVSS 0.112692f
C4166 IREF.n10 AVSS 0.112636f
C4167 IREF.t25 AVSS 0.120793f
C4168 IREF.n11 AVSS 0.16505f
C4169 IREF.n12 AVSS 0.061105f
C4170 IREF.n13 AVSS 0.235557f
C4171 IREF.n14 AVSS 0.235477f
C4172 IREF.t5 AVSS 0.120793f
C4173 IREF.n15 AVSS 0.16505f
C4174 IREF.n16 AVSS 0.060144f
C4175 IREF.n17 AVSS 0.112692f
C4176 IREF.n18 AVSS 0.112636f
C4177 IREF.t1 AVSS 0.239863f
C4178 IREF.n19 AVSS 0.390771f
C4179 IREF.t23 AVSS 0.25051f
C4180 IREF.t43 AVSS 0.046573f
C4181 IREF.t41 AVSS 0.046573f
C4182 IREF.n20 AVSS 0.188288f
C4183 IREF.n21 AVSS 0.63794f
C4184 IREF.t29 AVSS 0.186253f
C4185 IREF.n22 AVSS 0.543973f
C4186 IREF.t11 AVSS 0.186253f
C4187 IREF.n23 AVSS 0.536766f
C4188 IREF.n24 AVSS 0.120759f
C4189 IREF.t9 AVSS 0.242653f
C4190 IREF.t21 AVSS 0.046573f
C4191 IREF.t33 AVSS 0.046573f
C4192 IREF.n25 AVSS 0.118121f
C4193 IREF.n26 AVSS 0.185402f
C4194 IREF.n27 AVSS 0.392238f
C4195 IREF.n28 AVSS 0.594057f
C4196 IREF.n29 AVSS 0.0275f
C4197 IREF.t3 AVSS 0.046573f
C4198 IREF.t39 AVSS 0.046573f
C4199 IREF.n30 AVSS 0.117749f
C4200 IREF.t17 AVSS 0.046573f
C4201 IREF.t13 AVSS 0.046573f
C4202 IREF.n31 AVSS 0.107883f
C4203 IREF.n32 AVSS 0.635239f
C4204 IREF.n33 AVSS 0.594735f
C4205 IREF.t35 AVSS 0.122233f
C4206 IREF.n34 AVSS 0.16951f
C4207 IREF.t7 AVSS 0.113728f
C4208 IREF.n35 AVSS 0.194986f
C4209 IREF.n36 AVSS 0.373882f
C4210 IREF.n37 AVSS 3.57913f
C4211 IREF.n38 AVSS 2.71732f
C4212 IREF.n39 AVSS 2.76082f
C4213 IREF.n40 AVSS 0.096473f
C4214 IREF.n41 AVSS 0.0275f
C4215 IREF.n42 AVSS 0.0275f
C4216 IREF.n43 AVSS 0.16162f
C4217 IREF.n44 AVSS 0.049235f
C4218 IREF.t143 AVSS 0.388691f
C4219 IREF.n45 AVSS 0.307321f
C4220 IREF.n46 AVSS 0.0275f
C4221 IREF.n47 AVSS 0.147618f
C4222 IREF.n48 AVSS 0.0275f
C4223 IREF.n49 AVSS 0.064265f
C4224 IREF.n50 AVSS 0.050676f
C4225 IREF.n51 AVSS 0.177998f
C4226 IREF.t169 AVSS 0.388691f
C4227 IREF.n52 AVSS 0.187433f
C4228 IREF.n53 AVSS 0.049456f
C4229 IREF.t157 AVSS 0.388691f
C4230 IREF.n54 AVSS 0.187435f
C4231 IREF.n55 AVSS 0.049456f
C4232 IREF.n56 AVSS 0.058424f
C4233 IREF.n57 AVSS 0.062993f
C4234 IREF.t139 AVSS 0.388691f
C4235 IREF.n58 AVSS 0.187435f
C4236 IREF.n59 AVSS 0.073102f
C4237 IREF.n60 AVSS 0.063423f
C4238 IREF.n61 AVSS 0.049456f
C4239 IREF.n62 AVSS 0.173715f
C4240 IREF.n63 AVSS 0.162809f
C4241 IREF.n64 AVSS 0.049456f
C4242 IREF.n65 AVSS 0.0275f
C4243 IREF.n66 AVSS 0.059203f
C4244 IREF.n67 AVSS 0.0275f
C4245 IREF.n68 AVSS 0.050676f
C4246 IREF.n69 AVSS 0.050676f
C4247 IREF.n70 AVSS 0.162028f
C4248 IREF.n71 AVSS 0.050676f
C4249 IREF.n72 AVSS 0.0275f
C4250 IREF.n73 AVSS 0.042027f
C4251 IREF.n74 AVSS 0.042027f
C4252 IREF.n75 AVSS 0.147618f
C4253 IREF.n76 AVSS 0.042027f
C4254 IREF.n77 AVSS 0.042027f
C4255 IREF.n78 AVSS 0.0275f
C4256 IREF.n79 AVSS 0.057645f
C4257 IREF.t245 AVSS 0.388691f
C4258 IREF.n80 AVSS 0.187435f
C4259 IREF.n81 AVSS 0.070109f
C4260 IREF.n82 AVSS 0.088943f
C4261 IREF.n83 AVSS 0.093035f
C4262 IREF.n84 AVSS 0.058324f
C4263 IREF.n85 AVSS 0.16162f
C4264 IREF.n86 AVSS 0.163089f
C4265 IREF.t127 AVSS 0.388691f
C4266 IREF.n87 AVSS 0.184685f
C4267 IREF.n88 AVSS 0.047017f
C4268 IREF.n89 AVSS 0.0275f
C4269 IREF.n90 AVSS 0.049235f
C4270 IREF.n91 AVSS 0.049235f
C4271 IREF.n92 AVSS 0.163089f
C4272 IREF.n93 AVSS 0.047017f
C4273 IREF.t198 AVSS 0.388691f
C4274 IREF.n94 AVSS 0.260402f
C4275 IREF.n95 AVSS 0.083187f
C4276 IREF.n96 AVSS 0.082501f
C4277 IREF.n97 AVSS 0.0275f
C4278 IREF.n98 AVSS 0.049456f
C4279 IREF.n99 AVSS 0.162809f
C4280 IREF.n100 AVSS 0.050676f
C4281 IREF.t45 AVSS 0.388691f
C4282 IREF.n101 AVSS 0.187435f
C4283 IREF.n102 AVSS 0.049456f
C4284 IREF.n103 AVSS 0.0275f
C4285 IREF.n104 AVSS 0.050676f
C4286 IREF.n105 AVSS 0.050676f
C4287 IREF.t165 AVSS 0.388691f
C4288 IREF.n106 AVSS 0.187433f
C4289 IREF.n107 AVSS 0.042027f
C4290 IREF.n108 AVSS 0.0275f
C4291 IREF.n109 AVSS 0.042027f
C4292 IREF.n110 AVSS 0.042027f
C4293 IREF.n111 AVSS 0.057645f
C4294 IREF.n112 AVSS 0.311819f
C4295 IREF.t154 AVSS 0.388691f
C4296 IREF.n113 AVSS 0.187435f
C4297 IREF.n114 AVSS 0.0275f
C4298 IREF.n115 AVSS 0.0275f
C4299 IREF.n116 AVSS 0.173715f
C4300 IREF.n117 AVSS 0.0275f
C4301 IREF.n118 AVSS 0.049456f
C4302 IREF.n119 AVSS 0.049456f
C4303 IREF.n120 AVSS 0.0275f
C4304 IREF.n121 AVSS 0.050676f
C4305 IREF.n122 AVSS 0.162028f
C4306 IREF.n123 AVSS 0.042027f
C4307 IREF.t51 AVSS 0.388691f
C4308 IREF.n124 AVSS 0.187433f
C4309 IREF.n125 AVSS 0.050676f
C4310 IREF.n126 AVSS 0.0275f
C4311 IREF.n127 AVSS 0.042027f
C4312 IREF.n128 AVSS 0.042027f
C4313 IREF.n129 AVSS 0.057645f
C4314 IREF.n130 AVSS 0.876294f
C4315 IREF.n131 AVSS 0.096473f
C4316 IREF.n132 AVSS 0.0275f
C4317 IREF.n133 AVSS 0.0275f
C4318 IREF.n134 AVSS 0.16162f
C4319 IREF.n135 AVSS 0.049235f
C4320 IREF.t99 AVSS 0.388691f
C4321 IREF.n136 AVSS 0.307321f
C4322 IREF.n137 AVSS 0.0275f
C4323 IREF.n138 AVSS 0.147618f
C4324 IREF.n139 AVSS 0.0275f
C4325 IREF.n140 AVSS 0.064265f
C4326 IREF.n141 AVSS 0.050676f
C4327 IREF.n142 AVSS 0.177998f
C4328 IREF.t164 AVSS 0.388691f
C4329 IREF.n143 AVSS 0.187433f
C4330 IREF.n144 AVSS 0.049456f
C4331 IREF.t73 AVSS 0.388691f
C4332 IREF.n145 AVSS 0.187435f
C4333 IREF.n146 AVSS 0.049456f
C4334 IREF.n147 AVSS 0.058424f
C4335 IREF.n148 AVSS 0.311819f
C4336 IREF.n149 AVSS 0.0275f
C4337 IREF.n150 AVSS 0.147618f
C4338 IREF.n151 AVSS 0.0275f
C4339 IREF.n152 AVSS 0.064265f
C4340 IREF.n153 AVSS 0.050676f
C4341 IREF.n154 AVSS 0.177998f
C4342 IREF.t244 AVSS 0.388691f
C4343 IREF.n155 AVSS 0.187433f
C4344 IREF.n156 AVSS 0.049456f
C4345 IREF.t175 AVSS 0.388691f
C4346 IREF.n157 AVSS 0.187435f
C4347 IREF.n158 AVSS 0.049456f
C4348 IREF.n159 AVSS 0.058424f
C4349 IREF.n160 AVSS 0.094308f
C4350 IREF.n161 AVSS 0.0275f
C4351 IREF.n162 AVSS 0.038171f
C4352 IREF.n163 AVSS 0.0275f
C4353 IREF.n164 AVSS 0.171378f
C4354 IREF.n165 AVSS 0.049235f
C4355 IREF.t110 AVSS 0.388691f
C4356 IREF.n166 AVSS 0.317522f
C4357 IREF.n167 AVSS 0.0275f
C4358 IREF.n168 AVSS 0.048298f
C4359 IREF.n169 AVSS 0.049235f
C4360 IREF.n170 AVSS 0.116846f
C4361 IREF.n171 AVSS 0.050676f
C4362 IREF.n172 AVSS 0.048295f
C4363 IREF.n173 AVSS 0.049235f
C4364 IREF.n174 AVSS 0.048298f
C4365 IREF.n175 AVSS 0.049456f
C4366 IREF.n176 AVSS 0.048298f
C4367 IREF.n177 AVSS 0.103005f
C4368 IREF.n178 AVSS 0.048298f
C4369 IREF.n179 AVSS 0.098997f
C4370 IREF.t225 AVSS 0.388691f
C4371 IREF.n180 AVSS 0.186037f
C4372 IREF.n181 AVSS 0.04674f
C4373 IREF.n182 AVSS 0.063308f
C4374 IREF.n183 AVSS 0.049456f
C4375 IREF.n184 AVSS 0.124639f
C4376 IREF.n185 AVSS 0.125418f
C4377 IREF.n186 AVSS 0.049235f
C4378 IREF.n187 AVSS 0.0275f
C4379 IREF.n188 AVSS 0.037392f
C4380 IREF.t95 AVSS 0.388691f
C4381 IREF.n189 AVSS 0.151602f
C4382 IREF.n190 AVSS 0.04674f
C4383 IREF.n191 AVSS 0.0275f
C4384 IREF.n192 AVSS 0.050676f
C4385 IREF.n193 AVSS 0.124639f
C4386 IREF.n194 AVSS 0.129701f
C4387 IREF.n195 AVSS 0.049235f
C4388 IREF.n196 AVSS 0.0275f
C4389 IREF.n197 AVSS 0.032327f
C4390 IREF.t161 AVSS 0.388691f
C4391 IREF.n198 AVSS 0.156664f
C4392 IREF.n199 AVSS 0.048295f
C4393 IREF.n200 AVSS 0.046737f
C4394 IREF.n201 AVSS 0.0275f
C4395 IREF.n202 AVSS 0.042027f
C4396 IREF.n203 AVSS 0.042027f
C4397 IREF.n204 AVSS 0.10711f
C4398 IREF.n205 AVSS 0.048298f
C4399 IREF.n206 AVSS 0.049235f
C4400 IREF.n207 AVSS 0.0275f
C4401 IREF.n208 AVSS 0.009348f
C4402 IREF.t156 AVSS 0.388691f
C4403 IREF.n209 AVSS 0.179645f
C4404 IREF.n210 AVSS 0.084078f
C4405 IREF.n211 AVSS 0.088941f
C4406 IREF.n212 AVSS 0.093036f
C4407 IREF.n213 AVSS 0.058325f
C4408 IREF.n214 AVSS 0.171378f
C4409 IREF.n215 AVSS 0.172936f
C4410 IREF.t67 AVSS 0.388691f
C4411 IREF.n216 AVSS 0.187435f
C4412 IREF.n217 AVSS 0.049856f
C4413 IREF.n218 AVSS 0.0275f
C4414 IREF.n219 AVSS 0.049235f
C4415 IREF.n220 AVSS 0.049235f
C4416 IREF.n221 AVSS 0.172936f
C4417 IREF.n222 AVSS 0.049856f
C4418 IREF.t215 AVSS 0.388691f
C4419 IREF.n223 AVSS 0.267764f
C4420 IREF.n224 AVSS 0.083187f
C4421 IREF.n225 AVSS 0.049456f
C4422 IREF.t236 AVSS 0.388691f
C4423 IREF.n226 AVSS 0.150823f
C4424 IREF.n227 AVSS 0.124639f
C4425 IREF.n228 AVSS 0.0275f
C4426 IREF.n229 AVSS 0.037392f
C4427 IREF.n230 AVSS 0.050676f
C4428 IREF.t191 AVSS 0.388691f
C4429 IREF.n231 AVSS 0.151602f
C4430 IREF.n232 AVSS 0.124639f
C4431 IREF.n233 AVSS 0.0275f
C4432 IREF.n234 AVSS 0.032327f
C4433 IREF.n235 AVSS 0.042027f
C4434 IREF.t259 AVSS 0.388691f
C4435 IREF.n236 AVSS 0.156664f
C4436 IREF.n237 AVSS 0.116846f
C4437 IREF.n238 AVSS 0.0275f
C4438 IREF.n239 AVSS 0.10711f
C4439 IREF.n240 AVSS 0.009348f
C4440 IREF.n241 AVSS 0.042027f
C4441 IREF.n242 AVSS 0.311819f
C4442 IREF.t218 AVSS 0.388691f
C4443 IREF.n243 AVSS 0.179645f
C4444 IREF.n244 AVSS 0.0275f
C4445 IREF.n245 AVSS 0.048298f
C4446 IREF.n246 AVSS 0.049456f
C4447 IREF.n247 AVSS 0.048298f
C4448 IREF.n248 AVSS 0.049235f
C4449 IREF.n249 AVSS 0.049235f
C4450 IREF.n250 AVSS 0.048298f
C4451 IREF.n251 AVSS 0.050676f
C4452 IREF.n252 AVSS 0.048295f
C4453 IREF.n253 AVSS 0.049235f
C4454 IREF.n254 AVSS 0.048295f
C4455 IREF.n255 AVSS 0.042027f
C4456 IREF.n256 AVSS 0.048298f
C4457 IREF.n257 AVSS 0.094308f
C4458 IREF.n258 AVSS 0.0275f
C4459 IREF.n259 AVSS 0.058325f
C4460 IREF.n260 AVSS 0.049856f
C4461 IREF.n261 AVSS 0.049235f
C4462 IREF.t132 AVSS 0.388691f
C4463 IREF.n262 AVSS 0.187435f
C4464 IREF.t64 AVSS 0.388691f
C4465 IREF.n263 AVSS 0.267764f
C4466 IREF.n264 AVSS 0.0275f
C4467 IREF.n265 AVSS 0.217655f
C4468 IREF.t247 AVSS 0.388691f
C4469 IREF.n266 AVSS 0.150823f
C4470 IREF.n267 AVSS 0.049235f
C4471 IREF.n268 AVSS 0.04674f
C4472 IREF.n269 AVSS 0.125418f
C4473 IREF.n270 AVSS 0.0275f
C4474 IREF.t208 AVSS 0.388691f
C4475 IREF.n271 AVSS 0.151602f
C4476 IREF.n272 AVSS 0.049235f
C4477 IREF.n273 AVSS 0.04674f
C4478 IREF.n274 AVSS 0.129701f
C4479 IREF.n275 AVSS 0.0275f
C4480 IREF.t60 AVSS 0.388691f
C4481 IREF.n276 AVSS 0.156664f
C4482 IREF.n277 AVSS 0.049235f
C4483 IREF.n278 AVSS 0.046737f
C4484 IREF.n279 AVSS 0.10711f
C4485 IREF.n280 AVSS 0.091302f
C4486 IREF.n281 AVSS 0.048298f
C4487 IREF.t71 AVSS 0.388691f
C4488 IREF.n282 AVSS 0.179645f
C4489 IREF.n283 AVSS 0.061976f
C4490 IREF.n284 AVSS 0.009348f
C4491 IREF.n285 AVSS 0.048298f
C4492 IREF.n286 AVSS 0.100637f
C4493 IREF.n287 AVSS 0.042027f
C4494 IREF.n288 AVSS 0.042027f
C4495 IREF.n289 AVSS 0.116846f
C4496 IREF.n290 AVSS 0.048295f
C4497 IREF.n291 AVSS 0.049235f
C4498 IREF.n292 AVSS 0.0275f
C4499 IREF.n293 AVSS 0.032327f
C4500 IREF.n294 AVSS 0.048295f
C4501 IREF.n295 AVSS 0.050676f
C4502 IREF.n296 AVSS 0.050676f
C4503 IREF.n297 AVSS 0.124639f
C4504 IREF.n298 AVSS 0.048298f
C4505 IREF.n299 AVSS 0.049235f
C4506 IREF.n300 AVSS 0.0275f
C4507 IREF.n301 AVSS 0.037392f
C4508 IREF.n302 AVSS 0.048298f
C4509 IREF.n303 AVSS 0.049456f
C4510 IREF.n304 AVSS 0.049456f
C4511 IREF.n305 AVSS 0.124639f
C4512 IREF.n306 AVSS 0.048298f
C4513 IREF.n307 AVSS 0.049235f
C4514 IREF.n308 AVSS 0.0275f
C4515 IREF.n309 AVSS 0.038171f
C4516 IREF.n310 AVSS 0.091051f
C4517 IREF.n311 AVSS 0.082501f
C4518 IREF.n312 AVSS 0.083187f
C4519 IREF.n313 AVSS 0.0275f
C4520 IREF.n314 AVSS 0.049856f
C4521 IREF.n315 AVSS 0.172936f
C4522 IREF.n316 AVSS 0.171378f
C4523 IREF.n317 AVSS 0.049235f
C4524 IREF.n318 AVSS 0.0275f
C4525 IREF.n319 AVSS 0.049235f
C4526 IREF.n320 AVSS 0.172936f
C4527 IREF.n321 AVSS 0.171378f
C4528 IREF.t122 AVSS 0.388691f
C4529 IREF.n322 AVSS 0.317522f
C4530 IREF.n323 AVSS 0.093036f
C4531 IREF.n324 AVSS 0.088941f
C4532 IREF.n325 AVSS 0.084078f
C4533 IREF.t101 AVSS 0.388691f
C4534 IREF.n326 AVSS 0.179645f
C4535 IREF.n327 AVSS 0.009348f
C4536 IREF.n328 AVSS 0.0275f
C4537 IREF.n329 AVSS 0.049235f
C4538 IREF.n330 AVSS 0.048298f
C4539 IREF.n331 AVSS 0.10711f
C4540 IREF.n332 AVSS 0.116846f
C4541 IREF.n333 AVSS 0.042027f
C4542 IREF.n334 AVSS 0.0275f
C4543 IREF.n335 AVSS 0.046737f
C4544 IREF.t174 AVSS 0.388691f
C4545 IREF.n336 AVSS 0.156664f
C4546 IREF.n337 AVSS 0.032327f
C4547 IREF.n338 AVSS 0.0275f
C4548 IREF.n339 AVSS 0.049235f
C4549 IREF.n340 AVSS 0.129701f
C4550 IREF.n341 AVSS 0.124639f
C4551 IREF.n342 AVSS 0.050676f
C4552 IREF.n343 AVSS 0.0275f
C4553 IREF.n344 AVSS 0.04674f
C4554 IREF.t84 AVSS 0.388691f
C4555 IREF.n345 AVSS 0.151602f
C4556 IREF.n346 AVSS 0.037392f
C4557 IREF.n347 AVSS 0.0275f
C4558 IREF.n348 AVSS 0.049235f
C4559 IREF.n349 AVSS 0.125418f
C4560 IREF.n350 AVSS 0.124639f
C4561 IREF.n351 AVSS 0.049456f
C4562 IREF.n352 AVSS 0.0275f
C4563 IREF.n353 AVSS 0.04674f
C4564 IREF.t151 AVSS 0.388691f
C4565 IREF.n354 AVSS 0.150823f
C4566 IREF.n355 AVSS 0.038171f
C4567 IREF.n356 AVSS 0.091051f
C4568 IREF.n357 AVSS 0.306365f
C4569 IREF.n358 AVSS 0.306333f
C4570 IREF.n359 AVSS 0.087967f
C4571 IREF.n360 AVSS 0.311819f
C4572 IREF.n361 AVSS 0.0275f
C4573 IREF.n362 AVSS 0.048298f
C4574 IREF.n363 AVSS 0.048298f
C4575 IREF.n364 AVSS 0.049235f
C4576 IREF.n365 AVSS 0.049235f
C4577 IREF.n366 AVSS 0.048295f
C4578 IREF.n367 AVSS 0.046737f
C4579 IREF.n368 AVSS 0.0275f
C4580 IREF.n369 AVSS 0.050676f
C4581 IREF.n370 AVSS 0.048295f
C4582 IREF.n371 AVSS 0.129701f
C4583 IREF.n372 AVSS 0.049235f
C4584 IREF.n373 AVSS 0.049235f
C4585 IREF.n374 AVSS 0.048298f
C4586 IREF.n375 AVSS 0.04674f
C4587 IREF.n376 AVSS 0.0275f
C4588 IREF.n377 AVSS 0.049456f
C4589 IREF.n378 AVSS 0.048298f
C4590 IREF.n379 AVSS 0.125418f
C4591 IREF.n380 AVSS 0.049235f
C4592 IREF.n381 AVSS 0.049235f
C4593 IREF.n382 AVSS 0.048298f
C4594 IREF.n383 AVSS 0.04674f
C4595 IREF.n384 AVSS 0.0275f
C4596 IREF.n385 AVSS 0.082501f
C4597 IREF.n386 AVSS 0.091051f
C4598 IREF.n387 AVSS 0.217655f
C4599 IREF.n388 AVSS 0.876294f
C4600 IREF.n389 AVSS 4.31506f
C4601 IREF.n390 AVSS 0.289863f
C4602 IREF.n391 AVSS 0.0275f
C4603 IREF.n392 AVSS 0.16162f
C4604 IREF.n393 AVSS 0.049235f
C4605 IREF.t90 AVSS 0.388691f
C4606 IREF.n394 AVSS 0.307321f
C4607 IREF.n395 AVSS 0.0275f
C4608 IREF.t146 AVSS 0.388691f
C4609 IREF.n396 AVSS 0.187435f
C4610 IREF.n397 AVSS 0.042027f
C4611 IREF.n398 AVSS 0.147618f
C4612 IREF.n399 AVSS 0.050676f
C4613 IREF.t150 AVSS 0.388691f
C4614 IREF.n400 AVSS 0.187433f
C4615 IREF.n401 AVSS 0.050676f
C4616 IREF.n402 AVSS 0.059203f
C4617 IREF.n403 AVSS 0.049456f
C4618 IREF.n404 AVSS 0.173715f
C4619 IREF.t86 AVSS 0.388691f
C4620 IREF.n405 AVSS 0.187435f
C4621 IREF.n406 AVSS 0.073102f
C4622 IREF.t214 AVSS 0.388691f
C4623 IREF.n407 AVSS 0.187435f
C4624 IREF.n408 AVSS 0.062993f
C4625 IREF.n409 AVSS 0.058424f
C4626 IREF.n410 AVSS 0.063423f
C4627 IREF.n411 AVSS 0.049456f
C4628 IREF.n412 AVSS 0.0275f
C4629 IREF.n413 AVSS 0.049456f
C4630 IREF.n414 AVSS 0.162809f
C4631 IREF.n415 AVSS 0.049456f
C4632 IREF.n416 AVSS 0.0275f
C4633 IREF.n417 AVSS 0.050676f
C4634 IREF.n418 AVSS 0.177998f
C4635 IREF.n419 AVSS 0.162028f
C4636 IREF.n420 AVSS 0.050676f
C4637 IREF.n421 AVSS 0.042027f
C4638 IREF.n422 AVSS 0.0275f
C4639 IREF.n423 AVSS 0.064265f
C4640 IREF.n424 AVSS 0.0275f
C4641 IREF.n425 AVSS 0.042027f
C4642 IREF.n426 AVSS 0.042027f
C4643 IREF.n427 AVSS 0.147618f
C4644 IREF.n428 AVSS 0.057645f
C4645 IREF.n429 AVSS 0.0275f
C4646 IREF.n430 AVSS 0.096473f
C4647 IREF.n431 AVSS 0.070109f
C4648 IREF.n432 AVSS 0.088943f
C4649 IREF.n433 AVSS 0.093035f
C4650 IREF.n434 AVSS 0.058324f
C4651 IREF.n435 AVSS 0.16162f
C4652 IREF.n436 AVSS 0.163089f
C4653 IREF.t252 AVSS 0.388691f
C4654 IREF.n437 AVSS 0.184685f
C4655 IREF.n438 AVSS 0.047017f
C4656 IREF.n439 AVSS 0.0275f
C4657 IREF.n440 AVSS 0.049235f
C4658 IREF.n441 AVSS 0.049235f
C4659 IREF.n442 AVSS 0.163089f
C4660 IREF.n443 AVSS 0.047017f
C4661 IREF.t182 AVSS 0.388691f
C4662 IREF.n444 AVSS 0.260402f
C4663 IREF.n445 AVSS 0.083187f
C4664 IREF.n446 AVSS 0.0275f
C4665 IREF.n447 AVSS 0.082501f
C4666 IREF.t226 AVSS 0.388691f
C4667 IREF.n448 AVSS 0.187435f
C4668 IREF.n449 AVSS 0.070888f
C4669 IREF.n450 AVSS 0.22089f
C4670 IREF.n451 AVSS 0.0275f
C4671 IREF.n452 AVSS 0.049456f
C4672 IREF.n453 AVSS 0.173715f
C4673 IREF.n454 AVSS 0.162809f
C4674 IREF.n455 AVSS 0.049456f
C4675 IREF.n456 AVSS 0.0275f
C4676 IREF.n457 AVSS 0.059203f
C4677 IREF.n458 AVSS 0.0275f
C4678 IREF.n459 AVSS 0.050676f
C4679 IREF.n460 AVSS 0.050676f
C4680 IREF.n461 AVSS 0.162028f
C4681 IREF.n462 AVSS 0.050676f
C4682 IREF.n463 AVSS 0.0275f
C4683 IREF.n464 AVSS 0.042027f
C4684 IREF.n465 AVSS 0.042027f
C4685 IREF.n466 AVSS 0.147618f
C4686 IREF.n467 AVSS 0.042027f
C4687 IREF.n468 AVSS 0.042027f
C4688 IREF.n469 AVSS 0.0275f
C4689 IREF.n470 AVSS 0.057645f
C4690 IREF.t204 AVSS 0.388691f
C4691 IREF.n471 AVSS 0.187435f
C4692 IREF.n472 AVSS 0.070109f
C4693 IREF.n473 AVSS 0.311819f
C4694 IREF.n474 AVSS 0.0275f
C4695 IREF.n475 AVSS 0.311819f
C4696 IREF.t136 AVSS 0.388691f
C4697 IREF.n476 AVSS 0.187435f
C4698 IREF.n477 AVSS 0.070888f
C4699 IREF.n478 AVSS 0.311819f
C4700 IREF.n479 AVSS 0.0275f
C4701 IREF.n480 AVSS 0.049456f
C4702 IREF.n481 AVSS 0.173715f
C4703 IREF.n482 AVSS 0.162809f
C4704 IREF.n483 AVSS 0.049456f
C4705 IREF.n484 AVSS 0.0275f
C4706 IREF.n485 AVSS 0.059203f
C4707 IREF.n486 AVSS 0.0275f
C4708 IREF.n487 AVSS 0.050676f
C4709 IREF.n488 AVSS 0.050676f
C4710 IREF.n489 AVSS 0.162028f
C4711 IREF.n490 AVSS 0.050676f
C4712 IREF.n491 AVSS 0.0275f
C4713 IREF.n492 AVSS 0.042027f
C4714 IREF.n493 AVSS 0.042027f
C4715 IREF.n494 AVSS 0.147618f
C4716 IREF.n495 AVSS 0.042027f
C4717 IREF.n496 AVSS 0.042027f
C4718 IREF.n497 AVSS 0.0275f
C4719 IREF.n498 AVSS 0.057645f
C4720 IREF.t94 AVSS 0.388691f
C4721 IREF.n499 AVSS 0.187435f
C4722 IREF.n500 AVSS 0.070109f
C4723 IREF.n501 AVSS 0.088943f
C4724 IREF.n502 AVSS 0.093035f
C4725 IREF.n503 AVSS 0.058324f
C4726 IREF.n504 AVSS 0.16162f
C4727 IREF.n505 AVSS 0.163089f
C4728 IREF.t105 AVSS 0.388691f
C4729 IREF.n506 AVSS 0.184685f
C4730 IREF.n507 AVSS 0.047017f
C4731 IREF.n508 AVSS 0.0275f
C4732 IREF.n509 AVSS 0.049235f
C4733 IREF.n510 AVSS 0.049235f
C4734 IREF.n511 AVSS 0.163089f
C4735 IREF.n512 AVSS 0.047017f
C4736 IREF.t248 AVSS 0.388691f
C4737 IREF.n513 AVSS 0.260402f
C4738 IREF.n514 AVSS 0.083187f
C4739 IREF.n515 AVSS 0.082501f
C4740 IREF.n516 AVSS 0.0275f
C4741 IREF.n517 AVSS 0.049456f
C4742 IREF.n518 AVSS 0.162809f
C4743 IREF.n519 AVSS 0.050676f
C4744 IREF.t195 AVSS 0.388691f
C4745 IREF.n520 AVSS 0.187435f
C4746 IREF.n521 AVSS 0.049456f
C4747 IREF.n522 AVSS 0.0275f
C4748 IREF.n523 AVSS 0.050676f
C4749 IREF.n524 AVSS 0.050676f
C4750 IREF.t263 AVSS 0.388691f
C4751 IREF.n525 AVSS 0.187433f
C4752 IREF.n526 AVSS 0.042027f
C4753 IREF.n527 AVSS 0.0275f
C4754 IREF.n528 AVSS 0.042027f
C4755 IREF.n529 AVSS 0.042027f
C4756 IREF.n530 AVSS 0.057645f
C4757 IREF.t53 AVSS 0.388691f
C4758 IREF.n531 AVSS 0.187435f
C4759 IREF.n532 AVSS 0.100637f
C4760 IREF.n533 AVSS 0.073577f
C4761 IREF.n534 AVSS 0.06622f
C4762 IREF.n535 AVSS 0.042027f
C4763 IREF.n536 AVSS 0.147618f
C4764 IREF.n537 AVSS 0.147618f
C4765 IREF.n538 AVSS 0.064265f
C4766 IREF.n539 AVSS 0.0275f
C4767 IREF.n540 AVSS 0.050676f
C4768 IREF.n541 AVSS 0.162028f
C4769 IREF.n542 AVSS 0.177998f
C4770 IREF.n543 AVSS 0.059203f
C4771 IREF.n544 AVSS 0.0275f
C4772 IREF.n545 AVSS 0.049456f
C4773 IREF.n546 AVSS 0.049456f
C4774 IREF.n547 AVSS 0.173715f
C4775 IREF.n548 AVSS 0.058424f
C4776 IREF.t239 AVSS 0.388691f
C4777 IREF.n549 AVSS 0.187435f
C4778 IREF.n550 AVSS 0.070888f
C4779 IREF.n551 AVSS 0.22089f
C4780 IREF.n552 AVSS 0.289863f
C4781 IREF.n553 AVSS 4.31506f
C4782 IREF.n554 AVSS 0.094308f
C4783 IREF.n555 AVSS 0.0275f
C4784 IREF.n556 AVSS 0.038171f
C4785 IREF.n557 AVSS 0.0275f
C4786 IREF.n558 AVSS 0.171378f
C4787 IREF.n559 AVSS 0.049235f
C4788 IREF.t251 AVSS 0.388691f
C4789 IREF.n560 AVSS 0.317522f
C4790 IREF.n561 AVSS 0.0275f
C4791 IREF.n562 AVSS 0.048298f
C4792 IREF.n563 AVSS 0.049235f
C4793 IREF.n564 AVSS 0.116846f
C4794 IREF.n565 AVSS 0.050676f
C4795 IREF.n566 AVSS 0.048295f
C4796 IREF.n567 AVSS 0.049235f
C4797 IREF.n568 AVSS 0.048298f
C4798 IREF.n569 AVSS 0.049456f
C4799 IREF.n570 AVSS 0.048298f
C4800 IREF.n571 AVSS 0.049235f
C4801 IREF.n572 AVSS 0.048298f
C4802 IREF.n573 AVSS 0.311819f
C4803 IREF.n574 AVSS 0.091051f
C4804 IREF.n575 AVSS 0.0275f
C4805 IREF.t119 AVSS 0.388691f
C4806 IREF.n576 AVSS 0.179645f
C4807 IREF.n577 AVSS 0.042027f
C4808 IREF.n578 AVSS 0.10711f
C4809 IREF.n579 AVSS 0.0275f
C4810 IREF.n580 AVSS 0.046737f
C4811 IREF.n581 AVSS 0.050676f
C4812 IREF.n582 AVSS 0.124639f
C4813 IREF.n583 AVSS 0.0275f
C4814 IREF.t98 AVSS 0.388691f
C4815 IREF.n584 AVSS 0.151602f
C4816 IREF.n585 AVSS 0.049456f
C4817 IREF.n586 AVSS 0.124639f
C4818 IREF.n587 AVSS 0.0275f
C4819 IREF.t148 AVSS 0.388691f
C4820 IREF.n588 AVSS 0.150823f
C4821 IREF.n589 AVSS 0.083187f
C4822 IREF.n590 AVSS 0.0275f
C4823 IREF.t74 AVSS 0.388691f
C4824 IREF.n591 AVSS 0.179645f
C4825 IREF.n592 AVSS 0.042027f
C4826 IREF.n593 AVSS 0.10711f
C4827 IREF.n594 AVSS 0.0275f
C4828 IREF.n595 AVSS 0.046737f
C4829 IREF.n596 AVSS 0.050676f
C4830 IREF.n597 AVSS 0.124639f
C4831 IREF.n598 AVSS 0.0275f
C4832 IREF.t224 AVSS 0.388691f
C4833 IREF.n599 AVSS 0.151602f
C4834 IREF.n600 AVSS 0.049456f
C4835 IREF.n601 AVSS 0.124639f
C4836 IREF.n602 AVSS 0.098997f
C4837 IREF.t126 AVSS 0.388691f
C4838 IREF.n603 AVSS 0.186037f
C4839 IREF.n604 AVSS 0.063308f
C4840 IREF.n605 AVSS 0.04674f
C4841 IREF.n606 AVSS 0.048298f
C4842 IREF.n607 AVSS 0.103005f
C4843 IREF.n608 AVSS 0.049235f
C4844 IREF.n609 AVSS 0.125418f
C4845 IREF.n610 AVSS 0.037392f
C4846 IREF.n611 AVSS 0.048298f
C4847 IREF.n612 AVSS 0.049456f
C4848 IREF.n613 AVSS 0.0275f
C4849 IREF.n614 AVSS 0.04674f
C4850 IREF.n615 AVSS 0.048298f
C4851 IREF.n616 AVSS 0.049235f
C4852 IREF.n617 AVSS 0.049235f
C4853 IREF.n618 AVSS 0.129701f
C4854 IREF.t78 AVSS 0.388691f
C4855 IREF.n619 AVSS 0.156664f
C4856 IREF.n620 AVSS 0.032327f
C4857 IREF.n621 AVSS 0.048295f
C4858 IREF.n622 AVSS 0.050676f
C4859 IREF.n623 AVSS 0.0275f
C4860 IREF.n624 AVSS 0.042027f
C4861 IREF.n625 AVSS 0.116846f
C4862 IREF.n626 AVSS 0.048295f
C4863 IREF.n627 AVSS 0.049235f
C4864 IREF.n628 AVSS 0.049235f
C4865 IREF.n629 AVSS 0.048298f
C4866 IREF.n630 AVSS 0.009348f
C4867 IREF.n631 AVSS 0.048298f
C4868 IREF.n632 AVSS 0.0275f
C4869 IREF.n633 AVSS 0.058325f
C4870 IREF.n634 AVSS 0.049856f
C4871 IREF.n635 AVSS 0.049235f
C4872 IREF.t194 AVSS 0.388691f
C4873 IREF.n636 AVSS 0.187435f
C4874 IREF.t117 AVSS 0.388691f
C4875 IREF.n637 AVSS 0.267764f
C4876 IREF.n638 AVSS 0.0275f
C4877 IREF.n639 AVSS 0.049856f
C4878 IREF.n640 AVSS 0.172936f
C4879 IREF.n641 AVSS 0.171378f
C4880 IREF.n642 AVSS 0.049235f
C4881 IREF.n643 AVSS 0.0275f
C4882 IREF.n644 AVSS 0.049235f
C4883 IREF.n645 AVSS 0.172936f
C4884 IREF.n646 AVSS 0.171378f
C4885 IREF.t238 AVSS 0.388691f
C4886 IREF.n647 AVSS 0.317522f
C4887 IREF.n648 AVSS 0.093036f
C4888 IREF.n649 AVSS 0.088941f
C4889 IREF.n650 AVSS 0.084078f
C4890 IREF.n651 AVSS 0.094308f
C4891 IREF.n652 AVSS 0.284318f
C4892 IREF.n653 AVSS 0.217655f
C4893 IREF.n654 AVSS 0.038171f
C4894 IREF.n655 AVSS 0.091051f
C4895 IREF.n656 AVSS 0.082501f
C4896 IREF.n657 AVSS 0.0275f
C4897 IREF.n658 AVSS 0.04674f
C4898 IREF.n659 AVSS 0.048298f
C4899 IREF.n660 AVSS 0.049235f
C4900 IREF.n661 AVSS 0.049235f
C4901 IREF.n662 AVSS 0.125418f
C4902 IREF.n663 AVSS 0.037392f
C4903 IREF.n664 AVSS 0.048298f
C4904 IREF.n665 AVSS 0.049456f
C4905 IREF.n666 AVSS 0.0275f
C4906 IREF.n667 AVSS 0.04674f
C4907 IREF.n668 AVSS 0.048298f
C4908 IREF.n669 AVSS 0.049235f
C4909 IREF.n670 AVSS 0.049235f
C4910 IREF.n671 AVSS 0.129701f
C4911 IREF.t171 AVSS 0.388691f
C4912 IREF.n672 AVSS 0.156664f
C4913 IREF.n673 AVSS 0.032327f
C4914 IREF.n674 AVSS 0.048295f
C4915 IREF.n675 AVSS 0.050676f
C4916 IREF.n676 AVSS 0.0275f
C4917 IREF.n677 AVSS 0.042027f
C4918 IREF.n678 AVSS 0.116846f
C4919 IREF.n679 AVSS 0.048295f
C4920 IREF.n680 AVSS 0.049235f
C4921 IREF.n681 AVSS 0.049235f
C4922 IREF.n682 AVSS 0.048298f
C4923 IREF.n683 AVSS 0.009348f
C4924 IREF.n684 AVSS 0.048298f
C4925 IREF.n685 AVSS 0.0275f
C4926 IREF.n686 AVSS 0.311819f
C4927 IREF.n687 AVSS 0.087967f
C4928 IREF.n688 AVSS 0.306333f
C4929 IREF.n689 AVSS 0.306365f
C4930 IREF.n690 AVSS 0.0275f
C4931 IREF.n691 AVSS 0.038171f
C4932 IREF.t63 AVSS 0.388691f
C4933 IREF.n692 AVSS 0.150823f
C4934 IREF.n693 AVSS 0.04674f
C4935 IREF.n694 AVSS 0.0275f
C4936 IREF.n695 AVSS 0.049456f
C4937 IREF.n696 AVSS 0.124639f
C4938 IREF.n697 AVSS 0.125418f
C4939 IREF.n698 AVSS 0.049235f
C4940 IREF.n699 AVSS 0.0275f
C4941 IREF.n700 AVSS 0.037392f
C4942 IREF.t212 AVSS 0.388691f
C4943 IREF.n701 AVSS 0.151602f
C4944 IREF.n702 AVSS 0.04674f
C4945 IREF.n703 AVSS 0.0275f
C4946 IREF.n704 AVSS 0.050676f
C4947 IREF.n705 AVSS 0.124639f
C4948 IREF.n706 AVSS 0.129701f
C4949 IREF.n707 AVSS 0.049235f
C4950 IREF.n708 AVSS 0.0275f
C4951 IREF.n709 AVSS 0.032327f
C4952 IREF.t92 AVSS 0.388691f
C4953 IREF.n710 AVSS 0.156664f
C4954 IREF.n711 AVSS 0.048295f
C4955 IREF.n712 AVSS 0.046737f
C4956 IREF.n713 AVSS 0.0275f
C4957 IREF.n714 AVSS 0.042027f
C4958 IREF.n715 AVSS 0.042027f
C4959 IREF.n716 AVSS 0.10711f
C4960 IREF.n717 AVSS 0.048298f
C4961 IREF.n718 AVSS 0.049235f
C4962 IREF.n719 AVSS 0.0275f
C4963 IREF.n720 AVSS 0.009348f
C4964 IREF.t231 AVSS 0.388691f
C4965 IREF.n721 AVSS 0.179645f
C4966 IREF.n722 AVSS 0.084078f
C4967 IREF.n723 AVSS 0.088941f
C4968 IREF.n724 AVSS 0.093036f
C4969 IREF.n725 AVSS 0.058325f
C4970 IREF.n726 AVSS 0.171378f
C4971 IREF.n727 AVSS 0.172936f
C4972 IREF.t260 AVSS 0.388691f
C4973 IREF.n728 AVSS 0.187435f
C4974 IREF.n729 AVSS 0.049856f
C4975 IREF.n730 AVSS 0.0275f
C4976 IREF.n731 AVSS 0.049235f
C4977 IREF.n732 AVSS 0.049235f
C4978 IREF.n733 AVSS 0.172936f
C4979 IREF.n734 AVSS 0.049856f
C4980 IREF.t190 AVSS 0.388691f
C4981 IREF.n735 AVSS 0.267764f
C4982 IREF.n736 AVSS 0.083187f
C4983 IREF.n737 AVSS 0.049456f
C4984 IREF.t163 AVSS 0.388691f
C4985 IREF.n738 AVSS 0.150823f
C4986 IREF.n739 AVSS 0.124639f
C4987 IREF.n740 AVSS 0.0275f
C4988 IREF.n741 AVSS 0.037392f
C4989 IREF.n742 AVSS 0.050676f
C4990 IREF.t115 AVSS 0.388691f
C4991 IREF.n743 AVSS 0.151602f
C4992 IREF.n744 AVSS 0.124639f
C4993 IREF.n745 AVSS 0.0275f
C4994 IREF.n746 AVSS 0.032327f
C4995 IREF.n747 AVSS 0.042027f
C4996 IREF.t186 AVSS 0.388691f
C4997 IREF.n748 AVSS 0.156664f
C4998 IREF.n749 AVSS 0.116846f
C4999 IREF.n750 AVSS 0.061976f
C5000 IREF.n751 AVSS 0.10711f
C5001 IREF.n752 AVSS 0.009348f
C5002 IREF.n753 AVSS 0.042027f
C5003 IREF.t196 AVSS 0.388691f
C5004 IREF.n754 AVSS 0.179645f
C5005 IREF.n755 AVSS 0.091302f
C5006 IREF.n756 AVSS 0.100637f
C5007 IREF.n757 AVSS 0.048298f
C5008 IREF.n758 AVSS 0.048298f
C5009 IREF.n759 AVSS 0.049235f
C5010 IREF.n760 AVSS 0.049235f
C5011 IREF.n761 AVSS 0.048295f
C5012 IREF.n762 AVSS 0.046737f
C5013 IREF.n763 AVSS 0.0275f
C5014 IREF.n764 AVSS 0.050676f
C5015 IREF.n765 AVSS 0.048295f
C5016 IREF.n766 AVSS 0.129701f
C5017 IREF.n767 AVSS 0.049235f
C5018 IREF.n768 AVSS 0.049235f
C5019 IREF.n769 AVSS 0.048298f
C5020 IREF.n770 AVSS 0.04674f
C5021 IREF.n771 AVSS 0.0275f
C5022 IREF.n772 AVSS 0.049456f
C5023 IREF.n773 AVSS 0.048298f
C5024 IREF.n774 AVSS 0.125418f
C5025 IREF.n775 AVSS 0.049235f
C5026 IREF.n776 AVSS 0.049235f
C5027 IREF.n777 AVSS 0.048298f
C5028 IREF.n778 AVSS 0.04674f
C5029 IREF.n779 AVSS 0.0275f
C5030 IREF.n780 AVSS 0.082501f
C5031 IREF.n781 AVSS 0.091051f
C5032 IREF.n782 AVSS 0.217655f
C5033 IREF.n783 AVSS 0.284318f
C5034 IREF.n784 AVSS 2.76082f
C5035 IREF.n785 AVSS 2.76082f
C5036 IREF.n786 AVSS 0.227321f
C5037 IREF.n787 AVSS 0.0275f
C5038 IREF.n788 AVSS 0.046773f
C5039 IREF.n789 AVSS 0.0275f
C5040 IREF.n790 AVSS 0.046351f
C5041 IREF.n791 AVSS 0.049235f
C5042 IREF.t180 AVSS 0.388691f
C5043 IREF.n792 AVSS 0.186831f
C5044 IREF.n793 AVSS 0.0275f
C5045 IREF.n794 AVSS 0.046351f
C5046 IREF.n795 AVSS 0.049235f
C5047 IREF.t70 AVSS 0.388691f
C5048 IREF.n796 AVSS 0.152201f
C5049 IREF.n797 AVSS 0.049235f
C5050 IREF.t83 AVSS 0.388691f
C5051 IREF.n798 AVSS 0.152201f
C5052 IREF.n799 AVSS 0.084497f
C5053 IREF.t49 AVSS 0.388691f
C5054 IREF.n800 AVSS 0.152201f
C5055 IREF.n801 AVSS 0.049235f
C5056 IREF.t189 AVSS 0.388691f
C5057 IREF.n802 AVSS 0.152201f
C5058 IREF.n803 AVSS 0.049235f
C5059 IREF.t178 AVSS 0.388691f
C5060 IREF.n804 AVSS 0.202629f
C5061 IREF.t160 AVSS 0.397045f
C5062 IREF.n805 AVSS 0.28987f
C5063 IREF.n806 AVSS 0.178641f
C5064 IREF.n807 AVSS 0.046351f
C5065 IREF.n808 AVSS 0.046773f
C5066 IREF.n809 AVSS 0.013484f
C5067 IREF.n810 AVSS 0.0275f
C5068 IREF.n811 AVSS 0.049235f
C5069 IREF.n812 AVSS 0.046351f
C5070 IREF.n813 AVSS 0.046773f
C5071 IREF.n814 AVSS 0.013484f
C5072 IREF.n815 AVSS 0.0275f
C5073 IREF.n816 AVSS 1.04221f
C5074 IREF.n817 AVSS 0.227321f
C5075 IREF.n818 AVSS 0.0275f
C5076 IREF.n819 AVSS 0.046773f
C5077 IREF.n820 AVSS 0.0275f
C5078 IREF.n821 AVSS 0.046351f
C5079 IREF.t47 AVSS 0.388691f
C5080 IREF.n822 AVSS 0.202629f
C5081 IREF.t176 AVSS 0.397045f
C5082 IREF.n823 AVSS 0.28987f
C5083 IREF.n824 AVSS 0.178641f
C5084 IREF.n825 AVSS 0.049235f
C5085 IREF.n826 AVSS 0.046773f
C5086 IREF.n827 AVSS 0.013484f
C5087 IREF.t114 AVSS 0.388691f
C5088 IREF.n828 AVSS 0.152201f
C5089 IREF.n829 AVSS 0.046351f
C5090 IREF.n830 AVSS 0.049235f
C5091 IREF.n831 AVSS 0.049235f
C5092 IREF.n832 AVSS 0.0275f
C5093 IREF.n833 AVSS 0.013484f
C5094 IREF.t109 AVSS 0.388691f
C5095 IREF.n834 AVSS 0.152201f
C5096 IREF.n835 AVSS 0.130293f
C5097 IREF.t116 AVSS 0.388691f
C5098 IREF.n836 AVSS 0.314764f
C5099 IREF.t79 AVSS 0.388691f
C5100 IREF.n837 AVSS 0.258809f
C5101 IREF.t222 AVSS 0.388691f
C5102 IREF.n838 AVSS 0.313851f
C5103 IREF.n839 AVSS 0.046773f
C5104 IREF.n840 AVSS 0.049235f
C5105 IREF.n841 AVSS 0.013484f
C5106 IREF.n842 AVSS 0.049235f
C5107 IREF.t219 AVSS 0.388691f
C5108 IREF.n843 AVSS 0.152201f
C5109 IREF.t167 AVSS 0.388691f
C5110 IREF.n844 AVSS 0.172624f
C5111 IREF.n845 AVSS 0.058255f
C5112 IREF.n846 AVSS 0.013484f
C5113 IREF.n847 AVSS 0.049235f
C5114 IREF.t246 AVSS 0.388691f
C5115 IREF.n848 AVSS 0.152201f
C5116 IREF.t124 AVSS 0.388691f
C5117 IREF.n849 AVSS 0.152201f
C5118 IREF.n850 AVSS 0.049235f
C5119 IREF.t59 AVSS 0.388691f
C5120 IREF.n851 AVSS 0.152201f
C5121 IREF.n852 AVSS 0.229539f
C5122 IREF.n853 AVSS 0.0275f
C5123 IREF.n854 AVSS 0.039925f
C5124 IREF.n855 AVSS 0.0275f
C5125 IREF.n856 AVSS 0.048142f
C5126 IREF.n857 AVSS 0.049456f
C5127 IREF.n858 AVSS 0.015802f
C5128 IREF.n859 AVSS 0.0275f
C5129 IREF.n860 AVSS 0.039925f
C5130 IREF.n861 AVSS 0.050676f
C5131 IREF.n862 AVSS 0.016012f
C5132 IREF.n863 AVSS 0.049456f
C5133 IREF.t223 AVSS 0.388691f
C5134 IREF.n864 AVSS 0.152201f
C5135 IREF.t137 AVSS 0.388691f
C5136 IREF.n865 AVSS 0.152201f
C5137 IREF.n866 AVSS 0.042027f
C5138 IREF.n867 AVSS 0.017382f
C5139 IREF.n868 AVSS 0.050676f
C5140 IREF.t82 AVSS 0.388691f
C5141 IREF.n869 AVSS 0.192206f
C5142 IREF.t207 AVSS 0.39435f
C5143 IREF.n870 AVSS 0.271517f
C5144 IREF.n871 AVSS 0.151961f
C5145 IREF.n872 AVSS 0.016012f
C5146 IREF.n873 AVSS 0.048142f
C5147 IREF.t140 AVSS 0.388691f
C5148 IREF.n874 AVSS 0.152201f
C5149 IREF.n875 AVSS 0.043823f
C5150 IREF.n876 AVSS 0.050676f
C5151 IREF.n877 AVSS 0.0275f
C5152 IREF.n878 AVSS 0.042027f
C5153 IREF.n879 AVSS 0.039925f
C5154 IREF.n880 AVSS 0.039925f
C5155 IREF.n881 AVSS 0.015591f
C5156 IREF.n882 AVSS 0.0275f
C5157 IREF.n883 AVSS 0.229539f
C5158 IREF.n884 AVSS 0.130124f
C5159 IREF.t125 AVSS 0.388691f
C5160 IREF.n885 AVSS 0.31704f
C5161 IREF.t88 AVSS 0.388691f
C5162 IREF.n886 AVSS 0.258809f
C5163 IREF.t229 AVSS 0.388691f
C5164 IREF.n887 AVSS 0.317298f
C5165 IREF.n888 AVSS 0.130077f
C5166 IREF.n889 AVSS 0.087824f
C5167 IREF.n890 AVSS 0.0275f
C5168 IREF.n891 AVSS 0.015802f
C5169 IREF.n892 AVSS 0.046984f
C5170 IREF.t170 AVSS 0.388691f
C5171 IREF.n893 AVSS 0.152201f
C5172 IREF.n894 AVSS 0.044034f
C5173 IREF.n895 AVSS 0.049456f
C5174 IREF.n896 AVSS 0.0275f
C5175 IREF.n897 AVSS 0.050676f
C5176 IREF.n898 AVSS 0.048142f
C5177 IREF.n899 AVSS 0.043823f
C5178 IREF.t240 AVSS 0.388691f
C5179 IREF.n900 AVSS 0.152201f
C5180 IREF.n901 AVSS 0.017382f
C5181 IREF.n902 AVSS 0.0275f
C5182 IREF.n903 AVSS 0.042027f
C5183 IREF.n904 AVSS 0.042027f
C5184 IREF.n905 AVSS 0.039925f
C5185 IREF.n906 AVSS 0.015591f
C5186 IREF.t197 AVSS 0.388691f
C5187 IREF.n907 AVSS 0.174782f
C5188 IREF.n908 AVSS 0.312413f
C5189 IREF.t128 AVSS 0.388691f
C5190 IREF.n909 AVSS 0.170891f
C5191 IREF.n910 AVSS 0.312301f
C5192 IREF.n911 AVSS 0.0275f
C5193 IREF.n912 AVSS 0.049456f
C5194 IREF.n913 AVSS 0.046984f
C5195 IREF.n914 AVSS 0.044034f
C5196 IREF.t61 AVSS 0.388691f
C5197 IREF.n915 AVSS 0.152201f
C5198 IREF.n916 AVSS 0.016012f
C5199 IREF.n917 AVSS 0.0275f
C5200 IREF.n918 AVSS 0.050676f
C5201 IREF.n919 AVSS 0.050676f
C5202 IREF.n920 AVSS 0.043823f
C5203 IREF.t155 AVSS 0.388691f
C5204 IREF.n921 AVSS 0.152201f
C5205 IREF.n922 AVSS 0.017382f
C5206 IREF.n923 AVSS 0.039925f
C5207 IREF.n924 AVSS 0.042027f
C5208 IREF.n925 AVSS 0.042027f
C5209 IREF.n926 AVSS 0.0275f
C5210 IREF.n927 AVSS 0.015591f
C5211 IREF.t91 AVSS 0.388691f
C5212 IREF.n928 AVSS 0.152201f
C5213 IREF.n929 AVSS 0.130124f
C5214 IREF.t147 AVSS 0.388691f
C5215 IREF.n930 AVSS 0.31704f
C5216 IREF.t153 AVSS 0.388691f
C5217 IREF.n931 AVSS 0.258809f
C5218 IREF.t87 AVSS 0.388691f
C5219 IREF.n932 AVSS 0.317298f
C5220 IREF.n933 AVSS 0.044034f
C5221 IREF.n934 AVSS 0.050676f
C5222 IREF.t184 AVSS 0.388691f
C5223 IREF.n935 AVSS 0.152201f
C5224 IREF.t255 AVSS 0.388691f
C5225 IREF.n936 AVSS 0.195265f
C5226 IREF.t46 AVSS 0.396455f
C5227 IREF.n937 AVSS 0.289603f
C5228 IREF.n938 AVSS 0.177419f
C5229 IREF.n939 AVSS 0.043823f
C5230 IREF.n940 AVSS 0.048142f
C5231 IREF.n941 AVSS 0.016012f
C5232 IREF.n942 AVSS 0.0275f
C5233 IREF.n943 AVSS 0.049456f
C5234 IREF.n944 AVSS 0.049456f
C5235 IREF.n945 AVSS 0.046984f
C5236 IREF.n946 AVSS 0.015802f
C5237 IREF.t232 AVSS 0.388691f
C5238 IREF.n947 AVSS 0.152201f
C5239 IREF.n948 AVSS 0.130077f
C5240 IREF.n949 AVSS 0.087824f
C5241 IREF.n950 AVSS 1.04221f
C5242 IREF.n951 AVSS 4.1551f
C5243 IREF.n952 AVSS 0.284318f
C5244 IREF.n953 AVSS 0.013484f
C5245 IREF.n954 AVSS 0.049235f
C5246 IREF.t210 AVSS 0.388691f
C5247 IREF.n955 AVSS 0.152201f
C5248 IREF.t158 AVSS 0.388691f
C5249 IREF.n956 AVSS 0.152201f
C5250 IREF.n957 AVSS 0.049235f
C5251 IREF.t230 AVSS 0.388691f
C5252 IREF.n958 AVSS 0.190467f
C5253 IREF.t237 AVSS 0.393918f
C5254 IREF.n959 AVSS 0.274434f
C5255 IREF.n960 AVSS 0.150905f
C5256 IREF.n961 AVSS 0.013484f
C5257 IREF.n962 AVSS 0.046773f
C5258 IREF.n963 AVSS 0.046351f
C5259 IREF.n964 AVSS 0.049235f
C5260 IREF.n965 AVSS 0.0275f
C5261 IREF.n966 AVSS 0.013484f
C5262 IREF.n967 AVSS 0.046773f
C5263 IREF.n968 AVSS 0.046351f
C5264 IREF.n969 AVSS 0.049235f
C5265 IREF.n970 AVSS 0.0275f
C5266 IREF.n971 AVSS 0.084497f
C5267 IREF.n972 AVSS 0.129942f
C5268 IREF.t75 AVSS 0.388691f
C5269 IREF.n973 AVSS 0.313851f
C5270 IREF.t138 AVSS 0.388691f
C5271 IREF.n974 AVSS 0.258809f
C5272 IREF.t131 AVSS 0.388691f
C5273 IREF.n975 AVSS 0.314764f
C5274 IREF.n976 AVSS 0.130293f
C5275 IREF.n977 AVSS 0.227321f
C5276 IREF.n978 AVSS 0.0275f
C5277 IREF.n979 AVSS 0.013484f
C5278 IREF.n980 AVSS 0.046773f
C5279 IREF.n981 AVSS 0.046351f
C5280 IREF.n982 AVSS 0.049235f
C5281 IREF.n983 AVSS 0.0275f
C5282 IREF.n984 AVSS 0.013484f
C5283 IREF.n985 AVSS 0.046773f
C5284 IREF.n986 AVSS 0.046351f
C5285 IREF.n987 AVSS 0.049235f
C5286 IREF.n988 AVSS 0.0275f
C5287 IREF.n989 AVSS 0.049235f
C5288 IREF.n990 AVSS 0.046773f
C5289 IREF.n991 AVSS 0.046351f
C5290 IREF.t104 AVSS 0.388691f
C5291 IREF.n992 AVSS 0.186831f
C5292 IREF.n993 AVSS 0.318415f
C5293 IREF.n994 AVSS 0.314023f
C5294 IREF.n995 AVSS 0.0275f
C5295 IREF.n996 AVSS 0.013484f
C5296 IREF.n997 AVSS 0.046773f
C5297 IREF.n998 AVSS 0.046351f
C5298 IREF.n999 AVSS 0.049235f
C5299 IREF.n1000 AVSS 0.0275f
C5300 IREF.n1001 AVSS 0.049235f
C5301 IREF.n1002 AVSS 0.046773f
C5302 IREF.n1003 AVSS 0.046351f
C5303 IREF.t144 AVSS 0.388691f
C5304 IREF.n1004 AVSS 0.152201f
C5305 IREF.n1005 AVSS 0.013484f
C5306 IREF.n1006 AVSS 0.0275f
C5307 IREF.n1007 AVSS 0.049235f
C5308 IREF.n1008 AVSS 0.049235f
C5309 IREF.n1009 AVSS 0.046351f
C5310 IREF.t193 AVSS 0.388691f
C5311 IREF.n1010 AVSS 0.152201f
C5312 IREF.n1011 AVSS 0.013484f
C5313 IREF.n1012 AVSS 0.129942f
C5314 IREF.n1013 AVSS 0.084497f
C5315 IREF.n1014 AVSS 0.284318f
C5316 IREF.n1015 AVSS 4.1551f
C5317 IREF.n1016 AVSS 0.229539f
C5318 IREF.n1017 AVSS 0.0275f
C5319 IREF.n1018 AVSS 0.039925f
C5320 IREF.n1019 AVSS 0.0275f
C5321 IREF.n1020 AVSS 0.048142f
C5322 IREF.t111 AVSS 0.39435f
C5323 IREF.n1021 AVSS 0.271517f
C5324 IREF.t206 AVSS 0.388691f
C5325 IREF.n1022 AVSS 0.192206f
C5326 IREF.n1023 AVSS 0.016012f
C5327 IREF.n1024 AVSS 0.151961f
C5328 IREF.n1025 AVSS 0.050676f
C5329 IREF.n1026 AVSS 0.050676f
C5330 IREF.n1027 AVSS 0.043823f
C5331 IREF.t52 AVSS 0.388691f
C5332 IREF.n1028 AVSS 0.152201f
C5333 IREF.n1029 AVSS 0.017382f
C5334 IREF.n1030 AVSS 0.039925f
C5335 IREF.n1031 AVSS 0.042027f
C5336 IREF.n1032 AVSS 0.042027f
C5337 IREF.n1033 AVSS 0.0275f
C5338 IREF.n1034 AVSS 0.015591f
C5339 IREF.t48 AVSS 0.388691f
C5340 IREF.n1035 AVSS 0.152201f
C5341 IREF.n1036 AVSS 0.130124f
C5342 IREF.t256 AVSS 0.388691f
C5343 IREF.n1037 AVSS 0.31704f
C5344 IREF.t216 AVSS 0.388691f
C5345 IREF.n1038 AVSS 0.258809f
C5346 IREF.t135 AVSS 0.388691f
C5347 IREF.n1039 AVSS 0.317298f
C5348 IREF.n1040 AVSS 0.044034f
C5349 IREF.n1041 AVSS 0.050676f
C5350 IREF.t85 AVSS 0.388691f
C5351 IREF.n1042 AVSS 0.152201f
C5352 IREF.t152 AVSS 0.388691f
C5353 IREF.n1043 AVSS 0.152201f
C5354 IREF.n1044 AVSS 0.042027f
C5355 IREF.n1045 AVSS 0.015591f
C5356 IREF.n1046 AVSS 0.0275f
C5357 IREF.n1047 AVSS 0.044034f
C5358 IREF.n1048 AVSS 0.050676f
C5359 IREF.t188 AVSS 0.388691f
C5360 IREF.n1049 AVSS 0.152201f
C5361 IREF.t72 AVSS 0.388691f
C5362 IREF.n1050 AVSS 0.152201f
C5363 IREF.n1051 AVSS 0.042027f
C5364 IREF.n1052 AVSS 0.015591f
C5365 IREF.n1053 AVSS 0.289863f
C5366 IREF.t217 AVSS 0.388691f
C5367 IREF.n1054 AVSS 0.152201f
C5368 IREF.t142 AVSS 0.388691f
C5369 IREF.n1055 AVSS 0.152201f
C5370 IREF.n1056 AVSS 0.049456f
C5371 IREF.t96 AVSS 0.388691f
C5372 IREF.n1057 AVSS 0.152201f
C5373 IREF.n1058 AVSS 0.050676f
C5374 IREF.t166 AVSS 0.388691f
C5375 IREF.n1059 AVSS 0.195265f
C5376 IREF.t173 AVSS 0.396455f
C5377 IREF.n1060 AVSS 0.289603f
C5378 IREF.n1061 AVSS 0.177419f
C5379 IREF.n1062 AVSS 0.043823f
C5380 IREF.n1063 AVSS 0.048142f
C5381 IREF.n1064 AVSS 0.016012f
C5382 IREF.n1065 AVSS 0.0275f
C5383 IREF.n1066 AVSS 0.049456f
C5384 IREF.n1067 AVSS 0.044034f
C5385 IREF.n1068 AVSS 0.046984f
C5386 IREF.n1069 AVSS 0.015802f
C5387 IREF.n1070 AVSS 0.0275f
C5388 IREF.n1071 AVSS 0.087824f
C5389 IREF.n1072 AVSS 0.130077f
C5390 IREF.t213 AVSS 0.388691f
C5391 IREF.n1073 AVSS 0.317298f
C5392 IREF.t65 AVSS 0.388691f
C5393 IREF.n1074 AVSS 0.258809f
C5394 IREF.t56 AVSS 0.388691f
C5395 IREF.n1075 AVSS 0.31704f
C5396 IREF.n1076 AVSS 0.130124f
C5397 IREF.n1077 AVSS 0.229539f
C5398 IREF.n1078 AVSS 0.0275f
C5399 IREF.n1079 AVSS 0.042027f
C5400 IREF.n1080 AVSS 0.039925f
C5401 IREF.n1081 AVSS 0.039925f
C5402 IREF.n1082 AVSS 0.017382f
C5403 IREF.n1083 AVSS 0.0275f
C5404 IREF.n1084 AVSS 0.050676f
C5405 IREF.n1085 AVSS 0.043823f
C5406 IREF.n1086 AVSS 0.048142f
C5407 IREF.n1087 AVSS 0.016012f
C5408 IREF.n1088 AVSS 0.0275f
C5409 IREF.n1089 AVSS 0.049456f
C5410 IREF.n1090 AVSS 0.049456f
C5411 IREF.n1091 AVSS 0.046984f
C5412 IREF.n1092 AVSS 0.015802f
C5413 IREF.t258 AVSS 0.388691f
C5414 IREF.n1093 AVSS 0.170891f
C5415 IREF.n1094 AVSS 0.312301f
C5416 IREF.t102 AVSS 0.388691f
C5417 IREF.n1095 AVSS 0.174782f
C5418 IREF.n1096 AVSS 0.312413f
C5419 IREF.n1097 AVSS 0.0275f
C5420 IREF.n1098 AVSS 0.042027f
C5421 IREF.n1099 AVSS 0.039925f
C5422 IREF.n1100 AVSS 0.039925f
C5423 IREF.n1101 AVSS 0.017382f
C5424 IREF.n1102 AVSS 0.0275f
C5425 IREF.n1103 AVSS 0.050676f
C5426 IREF.n1104 AVSS 0.043823f
C5427 IREF.n1105 AVSS 0.048142f
C5428 IREF.n1106 AVSS 0.016012f
C5429 IREF.n1107 AVSS 0.0275f
C5430 IREF.n1108 AVSS 0.049456f
C5431 IREF.n1109 AVSS 0.049456f
C5432 IREF.n1110 AVSS 0.046984f
C5433 IREF.n1111 AVSS 0.015802f
C5434 IREF.t123 AVSS 0.388691f
C5435 IREF.n1112 AVSS 0.152201f
C5436 IREF.n1113 AVSS 0.130077f
C5437 IREF.n1114 AVSS 0.087824f
C5438 IREF.n1115 AVSS 0.289863f
C5439 IREF.n1116 AVSS 2.76082f
C5440 IREF.n1117 AVSS 2.5037f
C5441 IREF.n1118 AVSS 0.284318f
C5442 IREF.n1119 AVSS 0.227321f
C5443 IREF.n1120 AVSS 0.130293f
C5444 IREF.t120 AVSS 0.388691f
C5445 IREF.n1121 AVSS 0.314764f
C5446 IREF.t112 AVSS 0.388691f
C5447 IREF.n1122 AVSS 0.258809f
C5448 IREF.t177 AVSS 0.388691f
C5449 IREF.n1123 AVSS 0.313851f
C5450 IREF.n1124 AVSS 0.129942f
C5451 IREF.n1125 AVSS 0.013484f
C5452 IREF.n1126 AVSS 0.0275f
C5453 IREF.n1127 AVSS 0.049235f
C5454 IREF.n1128 AVSS 0.046351f
C5455 IREF.n1129 AVSS 0.046773f
C5456 IREF.n1130 AVSS 0.013484f
C5457 IREF.n1131 AVSS 0.0275f
C5458 IREF.n1132 AVSS 0.049235f
C5459 IREF.n1133 AVSS 0.046351f
C5460 IREF.n1134 AVSS 0.046773f
C5461 IREF.t183 AVSS 0.388691f
C5462 IREF.n1135 AVSS 0.152201f
C5463 IREF.n1136 AVSS 0.013484f
C5464 IREF.n1137 AVSS 0.0275f
C5465 IREF.n1138 AVSS 0.049235f
C5466 IREF.n1139 AVSS 0.049235f
C5467 IREF.n1140 AVSS 0.046773f
C5468 IREF.n1141 AVSS 0.013484f
C5469 IREF.t172 AVSS 0.388691f
C5470 IREF.n1142 AVSS 0.172624f
C5471 IREF.n1143 AVSS 0.314023f
C5472 IREF.n1144 AVSS 0.318415f
C5473 IREF.n1145 AVSS 0.058255f
C5474 IREF.n1146 AVSS 0.046351f
C5475 IREF.n1147 AVSS 0.046773f
C5476 IREF.t242 AVSS 0.388691f
C5477 IREF.n1148 AVSS 0.152201f
C5478 IREF.n1149 AVSS 0.013484f
C5479 IREF.n1150 AVSS 0.0275f
C5480 IREF.n1151 AVSS 0.049235f
C5481 IREF.n1152 AVSS 0.049235f
C5482 IREF.n1153 AVSS 0.046773f
C5483 IREF.n1154 AVSS 0.013484f
C5484 IREF.t77 AVSS 0.388691f
C5485 IREF.n1155 AVSS 0.152201f
C5486 IREF.n1156 AVSS 0.046351f
C5487 IREF.n1157 AVSS 0.049235f
C5488 IREF.n1158 AVSS 0.049235f
C5489 IREF.n1159 AVSS 0.0275f
C5490 IREF.n1160 AVSS 0.013484f
C5491 IREF.t129 AVSS 0.388691f
C5492 IREF.n1161 AVSS 0.152201f
C5493 IREF.n1162 AVSS 0.130293f
C5494 IREF.t262 AVSS 0.388691f
C5495 IREF.n1163 AVSS 0.314764f
C5496 IREF.t199 AVSS 0.388691f
C5497 IREF.n1164 AVSS 0.258809f
C5498 IREF.t257 AVSS 0.388691f
C5499 IREF.n1165 AVSS 0.313851f
C5500 IREF.n1166 AVSS 0.046773f
C5501 IREF.n1167 AVSS 0.049235f
C5502 IREF.n1168 AVSS 0.013484f
C5503 IREF.t254 AVSS 0.393918f
C5504 IREF.t103 AVSS 0.388691f
C5505 IREF.n1169 AVSS 0.190467f
C5506 IREF.n1170 AVSS 0.274434f
C5507 IREF.n1171 AVSS 0.150905f
C5508 IREF.n1172 AVSS 0.049235f
C5509 IREF.n1173 AVSS 0.046773f
C5510 IREF.n1174 AVSS 0.046351f
C5511 IREF.t209 AVSS 0.388691f
C5512 IREF.n1175 AVSS 0.152201f
C5513 IREF.n1176 AVSS 0.013484f
C5514 IREF.n1177 AVSS 0.0275f
C5515 IREF.n1178 AVSS 0.049235f
C5516 IREF.n1179 AVSS 0.049235f
C5517 IREF.n1180 AVSS 0.046351f
C5518 IREF.t221 AVSS 0.388691f
C5519 IREF.n1181 AVSS 0.152201f
C5520 IREF.n1182 AVSS 0.013484f
C5521 IREF.n1183 AVSS 0.129942f
C5522 IREF.n1184 AVSS 0.084497f
C5523 IREF.n1185 AVSS 0.284318f
C5524 IREF.n1186 AVSS 2.7547f
C5525 IREF.n1187 AVSS 3.42836f
C5526 IREF.n1188 AVSS 2.38166f
C5527 IREF.n1189 AVSS 0.289863f
C5528 IREF.t113 AVSS 0.388691f
C5529 IREF.n1190 AVSS 0.187435f
C5530 IREF.n1191 AVSS 0.0275f
C5531 IREF.n1192 AVSS 0.058324f
C5532 IREF.n1193 AVSS 0.047017f
C5533 IREF.n1194 AVSS 0.049235f
C5534 IREF.t220 AVSS 0.388691f
C5535 IREF.n1195 AVSS 0.184685f
C5536 IREF.t62 AVSS 0.388691f
C5537 IREF.n1196 AVSS 0.260402f
C5538 IREF.n1197 AVSS 0.0275f
C5539 IREF.t200 AVSS 0.388691f
C5540 IREF.n1198 AVSS 0.187435f
C5541 IREF.n1199 AVSS 0.049456f
C5542 IREF.n1200 AVSS 0.049456f
C5543 IREF.n1201 AVSS 0.049456f
C5544 IREF.t185 AVSS 0.388691f
C5545 IREF.n1202 AVSS 0.187435f
C5546 IREF.n1203 AVSS 0.050676f
C5547 IREF.n1204 AVSS 0.0275f
C5548 IREF.n1205 AVSS 0.050676f
C5549 IREF.n1206 AVSS 0.050676f
C5550 IREF.t93 AVSS 0.388691f
C5551 IREF.n1207 AVSS 0.187433f
C5552 IREF.n1208 AVSS 0.042027f
C5553 IREF.n1209 AVSS 0.0275f
C5554 IREF.n1210 AVSS 0.042027f
C5555 IREF.n1211 AVSS 0.042027f
C5556 IREF.n1212 AVSS 0.057645f
C5557 IREF.t235 AVSS 0.388691f
C5558 IREF.n1213 AVSS 0.187435f
C5559 IREF.n1214 AVSS 0.100637f
C5560 IREF.n1215 AVSS 0.073577f
C5561 IREF.n1216 AVSS 0.06622f
C5562 IREF.n1217 AVSS 0.042027f
C5563 IREF.n1218 AVSS 0.147618f
C5564 IREF.n1219 AVSS 0.147618f
C5565 IREF.n1220 AVSS 0.064265f
C5566 IREF.n1221 AVSS 0.0275f
C5567 IREF.n1222 AVSS 0.050676f
C5568 IREF.n1223 AVSS 0.162028f
C5569 IREF.n1224 AVSS 0.177998f
C5570 IREF.n1225 AVSS 0.059203f
C5571 IREF.n1226 AVSS 0.0275f
C5572 IREF.n1227 AVSS 0.049456f
C5573 IREF.n1228 AVSS 0.162809f
C5574 IREF.n1229 AVSS 0.173715f
C5575 IREF.n1230 AVSS 0.058424f
C5576 IREF.n1231 AVSS 0.0275f
C5577 IREF.n1232 AVSS 0.22089f
C5578 IREF.n1233 AVSS 0.070888f
C5579 IREF.n1234 AVSS 0.082501f
C5580 IREF.n1235 AVSS 0.083187f
C5581 IREF.n1236 AVSS 0.0275f
C5582 IREF.n1237 AVSS 0.047017f
C5583 IREF.n1238 AVSS 0.163089f
C5584 IREF.n1239 AVSS 0.16162f
C5585 IREF.n1240 AVSS 0.049235f
C5586 IREF.n1241 AVSS 0.0275f
C5587 IREF.n1242 AVSS 0.049235f
C5588 IREF.n1243 AVSS 0.163089f
C5589 IREF.n1244 AVSS 0.16162f
C5590 IREF.t69 AVSS 0.388691f
C5591 IREF.n1245 AVSS 0.307321f
C5592 IREF.n1246 AVSS 0.093035f
C5593 IREF.n1247 AVSS 0.088943f
C5594 IREF.n1248 AVSS 0.070109f
C5595 IREF.n1249 AVSS 0.096473f
C5596 IREF.n1250 AVSS 0.0275f
C5597 IREF.n1251 AVSS 0.042027f
C5598 IREF.n1252 AVSS 0.147618f
C5599 IREF.n1253 AVSS 0.147618f
C5600 IREF.n1254 AVSS 0.064265f
C5601 IREF.n1255 AVSS 0.0275f
C5602 IREF.n1256 AVSS 0.050676f
C5603 IREF.n1257 AVSS 0.050676f
C5604 IREF.n1258 AVSS 0.177998f
C5605 IREF.n1259 AVSS 0.059203f
C5606 IREF.t227 AVSS 0.388691f
C5607 IREF.n1260 AVSS 0.187435f
C5608 IREF.n1261 AVSS 0.162809f
C5609 IREF.n1262 AVSS 0.049456f
C5610 IREF.n1263 AVSS 0.049456f
C5611 IREF.n1264 AVSS 0.0275f
C5612 IREF.n1265 AVSS 0.058424f
C5613 IREF.t162 AVSS 0.388691f
C5614 IREF.n1266 AVSS 0.187435f
C5615 IREF.n1267 AVSS 0.070888f
C5616 IREF.n1268 AVSS 0.311819f
C5617 IREF.n1269 AVSS 0.311819f
C5618 IREF.n1270 AVSS 0.070109f
C5619 IREF.n1271 AVSS 0.311819f
C5620 IREF.n1272 AVSS 0.0275f
C5621 IREF.n1273 AVSS 0.042027f
C5622 IREF.n1274 AVSS 0.147618f
C5623 IREF.n1275 AVSS 0.147618f
C5624 IREF.n1276 AVSS 0.064265f
C5625 IREF.n1277 AVSS 0.0275f
C5626 IREF.n1278 AVSS 0.050676f
C5627 IREF.n1279 AVSS 0.162028f
C5628 IREF.n1280 AVSS 0.177998f
C5629 IREF.n1281 AVSS 0.059203f
C5630 IREF.n1282 AVSS 0.0275f
C5631 IREF.n1283 AVSS 0.049456f
C5632 IREF.n1284 AVSS 0.049456f
C5633 IREF.n1285 AVSS 0.173715f
C5634 IREF.n1286 AVSS 0.058424f
C5635 IREF.t58 AVSS 0.388691f
C5636 IREF.n1287 AVSS 0.187435f
C5637 IREF.n1288 AVSS 0.070888f
C5638 IREF.n1289 AVSS 0.22089f
C5639 IREF.n1290 AVSS 0.289863f
C5640 IREF.n1291 AVSS 2.38166f
C5641 IREF.n1292 AVSS 16.601f
C5642 IREF.t22 AVSS 0.438216f
C5643 IREF.t42 AVSS 0.420591f
C5644 IREF.n1293 AVSS 0.569166f
C5645 IREF.t40 AVSS 0.420597f
C5646 IREF.n1294 AVSS 0.302623f
C5647 IREF.t28 AVSS 0.420597f
C5648 IREF.n1295 AVSS 0.33055f
C5649 IREF.t211 AVSS 0.420706f
C5650 IREF.n1296 AVSS 0.332558f
C5651 IREF.t241 AVSS 0.420597f
C5652 IREF.n1297 AVSS 0.304744f
C5653 IREF.t249 AVSS 0.420603f
C5654 IREF.n1298 AVSS 0.259935f
C5655 IREF.t8 AVSS 0.438425f
C5656 IREF.t32 AVSS 0.420574f
C5657 IREF.n1299 AVSS 0.57299f
C5658 IREF.t20 AVSS 0.420574f
C5659 IREF.n1300 AVSS 0.302752f
C5660 IREF.t10 AVSS 0.420574f
C5661 IREF.n1301 AVSS 0.306188f
C5662 IREF.n1302 AVSS 0.178333f
C5663 IREF.t50 AVSS 0.438216f
C5664 IREF.t187 AVSS 0.420591f
C5665 IREF.n1303 AVSS 0.569166f
C5666 IREF.t201 AVSS 0.420597f
C5667 IREF.n1304 AVSS 0.302623f
C5668 IREF.t233 AVSS 0.420597f
C5669 IREF.n1305 AVSS 0.33055f
C5670 IREF.t118 AVSS 0.420706f
C5671 IREF.n1306 AVSS 0.332558f
C5672 IREF.t159 AVSS 0.420597f
C5673 IREF.n1307 AVSS 0.304744f
C5674 IREF.t168 AVSS 0.420603f
C5675 IREF.n1308 AVSS 0.259935f
C5676 IREF.t141 AVSS 0.438425f
C5677 IREF.t228 AVSS 0.420574f
C5678 IREF.n1309 AVSS 0.57299f
C5679 IREF.t76 AVSS 0.420574f
C5680 IREF.n1310 AVSS 0.302752f
C5681 IREF.t130 AVSS 0.420574f
C5682 IREF.n1311 AVSS 0.306188f
C5683 IREF.n1312 AVSS 0.100181f
C5684 IREF.n1313 AVSS 1.55438f
C5685 IREF.t179 AVSS 0.441063f
C5686 IREF.t97 AVSS 0.420591f
C5687 IREF.n1314 AVSS 0.612228f
C5688 IREF.t107 AVSS 0.420597f
C5689 IREF.n1315 AVSS 0.302623f
C5690 IREF.t145 AVSS 0.420597f
C5691 IREF.n1316 AVSS 0.33055f
C5692 IREF.t2 AVSS 0.420706f
C5693 IREF.n1317 AVSS 0.332558f
C5694 IREF.t38 AVSS 0.420597f
C5695 IREF.n1318 AVSS 0.304744f
C5696 IREF.t34 AVSS 0.420603f
C5697 IREF.n1319 AVSS 0.259935f
C5698 IREF.t55 AVSS 0.438686f
C5699 IREF.t133 AVSS 0.420574f
C5700 IREF.n1320 AVSS 0.576943f
C5701 IREF.t202 AVSS 0.420574f
C5702 IREF.n1321 AVSS 0.302752f
C5703 IREF.t261 AVSS 0.420574f
C5704 IREF.n1322 AVSS 0.306188f
C5705 IREF.n1323 AVSS 0.100181f
C5706 IREF.n1324 AVSS 1.03598f
C5707 IREF.t106 AVSS 0.438423f
C5708 IREF.t243 AVSS 0.420591f
C5709 IREF.n1325 AVSS 0.572286f
C5710 IREF.t253 AVSS 0.420597f
C5711 IREF.n1326 AVSS 0.302623f
C5712 IREF.t81 AVSS 0.420597f
C5713 IREF.n1327 AVSS 0.33055f
C5714 IREF.t16 AVSS 0.420706f
C5715 IREF.n1328 AVSS 0.332558f
C5716 IREF.t12 AVSS 0.420597f
C5717 IREF.n1329 AVSS 0.304744f
C5718 IREF.t6 AVSS 0.420603f
C5719 IREF.n1330 AVSS 0.259935f
C5720 IREF.t203 AVSS 0.438219f
C5721 IREF.t66 AVSS 0.420574f
C5722 IREF.n1331 AVSS 0.56987f
C5723 IREF.t121 AVSS 0.420574f
C5724 IREF.n1332 AVSS 0.302752f
C5725 IREF.t192 AVSS 0.420574f
C5726 IREF.n1333 AVSS 0.306188f
C5727 IREF.n1334 AVSS 0.100181f
C5728 IREF.n1335 AVSS 1.04418f
C5729 IREF.t181 AVSS 0.438216f
C5730 IREF.t100 AVSS 0.420591f
C5731 IREF.n1336 AVSS 0.569166f
C5732 IREF.t108 AVSS 0.420597f
C5733 IREF.n1337 AVSS 0.302623f
C5734 IREF.t149 AVSS 0.420597f
C5735 IREF.n1338 AVSS 0.33055f
C5736 IREF.t250 AVSS 0.420706f
C5737 IREF.n1339 AVSS 0.332558f
C5738 IREF.t80 AVSS 0.420597f
C5739 IREF.n1340 AVSS 0.304744f
C5740 IREF.t89 AVSS 0.420603f
C5741 IREF.n1341 AVSS 0.259935f
C5742 IREF.t57 AVSS 0.438425f
C5743 IREF.t134 AVSS 0.420574f
C5744 IREF.n1342 AVSS 0.57299f
C5745 IREF.t205 AVSS 0.420574f
C5746 IREF.n1343 AVSS 0.302752f
C5747 IREF.t44 AVSS 0.420574f
C5748 IREF.n1344 AVSS 0.306188f
C5749 IREF.n1345 AVSS 0.100181f
C5750 IREF.n1346 AVSS 0.576454f
C5751 IREF.n1347 AVSS 0.0275f
C5752 IREF.n1348 AVSS 0.046351f
C5753 IREF.n1349 AVSS 0.049124f
C5754 IREF.t36 AVSS 0.388691f
C5755 IREF.n1350 AVSS 0.202806f
C5756 IREF.t18 AVSS 0.397064f
C5757 IREF.n1351 AVSS 0.289887f
C5758 IREF.n1352 AVSS 0.178643f
C5759 IREF.n1353 AVSS 0.046351f
C5760 IREF.n1354 AVSS 0.046667f
C5761 IREF.t30 AVSS 0.388691f
C5762 IREF.n1355 AVSS 0.152201f
C5763 IREF.n1356 AVSS 0.013484f
C5764 IREF.n1357 AVSS 0.0275f
C5765 IREF.n1358 AVSS 0.049235f
C5766 IREF.n1359 AVSS 0.049235f
C5767 IREF.n1360 AVSS 0.046773f
C5768 IREF.n1361 AVSS 0.013484f
C5769 IREF.t24 AVSS 0.388691f
C5770 IREF.n1362 AVSS 0.177935f
C5771 IREF.n1363 AVSS 0.093106f
C5772 IREF.t234 AVSS 0.420706f
C5773 IREF.n1364 AVSS 0.317388f
C5774 IREF.t54 AVSS 0.420597f
C5775 IREF.n1365 AVSS 0.304744f
C5776 IREF.t68 AVSS 0.420603f
C5777 IREF.n1366 AVSS 0.259935f
C5778 IREF.t4 AVSS 0.388691f
C5779 IREF.n1367 AVSS 0.187503f
C5780 IREF.n1368 AVSS 0.049235f
C5781 IREF.t14 AVSS 0.388691f
C5782 IREF.n1369 AVSS 0.046773f
C5783 IREF.t0 AVSS 0.397119f
C5784 IREF.n1370 AVSS 0.290198f
C5785 IREF.t26 AVSS 0.388691f
C5786 IREF.n1371 AVSS 0.203244f
C5787 IREF.n1372 AVSS 0.046773f
C5788 IREF.n1373 AVSS 0.180994f
C5789 IREF.n1374 AVSS 0.049235f
C5790 IREF.n1375 AVSS 0.0275f
C5791 IREF.n1376 AVSS 0.165263f
C5792 IREF.n1377 AVSS 0.046773f
C5793 IREF.n1378 AVSS 0.046773f
C5794 IREF.n1379 AVSS 0.058255f
C5795 IREF.n1380 AVSS 0.079507f
C5796 IREF.n1381 AVSS 0.092525f
C5797 IREF.n1382 AVSS 1.60249f
C5798 IREF.n1383 AVSS 14.0357f
C5799 IREF.n1384 AVSS 2.45472f
C5800 IREF.n1385 AVSS 0.01375f
C5801 IREF.n1386 AVSS 0.014194f
C5802 IREF.n1387 AVSS 0.007374f
C5803 a_5396_8177.n0 AVSS 1.20526f
C5804 a_5396_8177.n1 AVSS 1.04691f
C5805 a_5396_8177.n2 AVSS 1.14821f
C5806 a_5396_8177.n3 AVSS 1.16512f
C5807 a_5396_8177.n4 AVSS 1.16506f
C5808 a_5396_8177.n5 AVSS 0.618667f
C5809 a_5396_8177.n6 AVSS 1.04691f
C5810 a_5396_8177.n7 AVSS 1.14827f
C5811 a_5396_8177.n8 AVSS 1.36794f
C5812 a_5396_8177.n9 AVSS 1.20526f
C5813 a_5396_8177.n10 AVSS 1.04691f
C5814 a_5396_8177.n11 AVSS 1.14827f
C5815 a_5396_8177.n12 AVSS 0.784419f
C5816 a_5396_8177.n13 AVSS 1.16507f
C5817 a_5396_8177.n14 AVSS 1.16506f
C5818 a_5396_8177.n15 AVSS 0.618667f
C5819 a_5396_8177.n16 AVSS 1.04691f
C5820 a_5396_8177.n17 AVSS 1.14827f
C5821 a_5396_8177.n18 AVSS 1.36794f
C5822 a_5396_8177.n19 AVSS 0.756645f
C5823 a_5396_8177.n20 AVSS 1.21829f
C5824 a_5396_8177.n21 AVSS 1.21828f
C5825 a_5396_8177.n22 AVSS 1.18637f
C5826 a_5396_8177.n23 AVSS 0.489163f
C5827 a_5396_8177.n24 AVSS 1.21829f
C5828 a_5396_8177.n25 AVSS 1.71656f
C5829 a_5396_8177.n26 AVSS 1.52625f
C5830 a_5396_8177.n27 AVSS 1.21829f
C5831 a_5396_8177.n28 AVSS 1.21828f
C5832 a_5396_8177.n29 AVSS 1.18637f
C5833 a_5396_8177.n30 AVSS 0.489163f
C5834 a_5396_8177.n31 AVSS 1.21829f
C5835 a_5396_8177.n32 AVSS 1.71656f
C5836 a_5396_8177.n33 AVSS 0.784419f
C5837 a_5396_8177.t51 AVSS 0.095293f
C5838 a_5396_8177.t32 AVSS 0.403593f
C5839 a_5396_8177.t73 AVSS 0.40307f
C5840 a_5396_8177.t44 AVSS 0.095293f
C5841 a_5396_8177.t25 AVSS 0.095293f
C5842 a_5396_8177.n34 AVSS 0.411692f
C5843 a_5396_8177.t53 AVSS 0.539266f
C5844 a_5396_8177.n35 AVSS 6.06825f
C5845 a_5396_8177.n36 AVSS 4.50976f
C5846 a_5396_8177.t38 AVSS 0.533524f
C5847 a_5396_8177.t18 AVSS 0.095293f
C5848 a_5396_8177.t84 AVSS 0.095293f
C5849 a_5396_8177.n37 AVSS 0.41253f
C5850 a_5396_8177.n38 AVSS 1.35792f
C5851 a_5396_8177.t66 AVSS 0.404415f
C5852 a_5396_8177.n39 AVSS 1.14932f
C5853 a_5396_8177.t2 AVSS 0.400953f
C5854 a_5396_8177.n40 AVSS 1.04137f
C5855 a_5396_8177.t0 AVSS 0.533524f
C5856 a_5396_8177.t68 AVSS 0.095293f
C5857 a_5396_8177.t47 AVSS 0.095293f
C5858 a_5396_8177.n41 AVSS 0.41253f
C5859 a_5396_8177.n42 AVSS 1.35792f
C5860 a_5396_8177.t28 AVSS 0.404415f
C5861 a_5396_8177.n43 AVSS 1.14932f
C5862 a_5396_8177.t52 AVSS 0.400953f
C5863 a_5396_8177.n44 AVSS 1.04137f
C5864 a_5396_8177.t41 AVSS 0.541038f
C5865 a_5396_8177.t33 AVSS 0.095293f
C5866 a_5396_8177.t14 AVSS 0.095293f
C5867 a_5396_8177.n45 AVSS 0.41253f
C5868 a_5396_8177.n46 AVSS 1.21102f
C5869 a_5396_8177.n47 AVSS 0.928418f
C5870 a_5396_8177.t61 AVSS 0.400953f
C5871 a_5396_8177.n48 AVSS 1.04137f
C5872 a_5396_8177.t21 AVSS 0.404415f
C5873 a_5396_8177.n49 AVSS 1.14932f
C5874 a_5396_8177.t76 AVSS 0.095293f
C5875 a_5396_8177.t40 AVSS 0.095293f
C5876 a_5396_8177.n50 AVSS 0.41253f
C5877 a_5396_8177.n51 AVSS 0.78412f
C5878 a_5396_8177.t6 AVSS 0.400953f
C5879 a_5396_8177.n52 AVSS 1.15658f
C5880 a_5396_8177.t54 AVSS 0.404302f
C5881 a_5396_8177.n53 AVSS 1.16606f
C5882 a_5396_8177.t22 AVSS 0.095293f
C5883 a_5396_8177.t85 AVSS 0.095293f
C5884 a_5396_8177.n54 AVSS 0.41253f
C5885 a_5396_8177.n55 AVSS 0.619074f
C5886 a_5396_8177.n56 AVSS 0.928418f
C5887 a_5396_8177.t24 AVSS 0.234869f
C5888 a_5396_8177.t29 AVSS 0.28657f
C5889 a_5396_8177.n57 AVSS 1.53577f
C5890 a_5396_8177.t83 AVSS 0.095293f
C5891 a_5396_8177.t63 AVSS 0.095293f
C5892 a_5396_8177.n58 AVSS 0.22302f
C5893 a_5396_8177.t1 AVSS 0.095293f
C5894 a_5396_8177.t69 AVSS 0.095293f
C5895 a_5396_8177.n59 AVSS 0.283728f
C5896 a_5396_8177.n60 AVSS 0.645783f
C5897 a_5396_8177.n61 AVSS 1.41165f
C5898 a_5396_8177.t72 AVSS 0.095293f
C5899 a_5396_8177.t50 AVSS 0.095293f
C5900 a_5396_8177.n62 AVSS 0.22302f
C5901 a_5396_8177.t74 AVSS 0.095293f
C5902 a_5396_8177.t55 AVSS 0.095293f
C5903 a_5396_8177.n63 AVSS 0.283728f
C5904 a_5396_8177.n64 AVSS 0.645783f
C5905 a_5396_8177.n65 AVSS 1.12242f
C5906 a_5396_8177.t12 AVSS 0.234869f
C5907 a_5396_8177.t17 AVSS 0.28657f
C5908 a_5396_8177.n66 AVSS 0.839828f
C5909 a_5396_8177.n67 AVSS 1.71657f
C5910 a_5396_8177.n68 AVSS 1.80896f
C5911 a_5396_8177.n69 AVSS 5.47384f
C5912 a_5396_8177.t11 AVSS 0.538544f
C5913 a_5396_8177.t81 AVSS 0.095293f
C5914 a_5396_8177.t58 AVSS 0.095293f
C5915 a_5396_8177.n70 AVSS 0.411692f
C5916 a_5396_8177.t39 AVSS 0.403593f
C5917 a_5396_8177.t64 AVSS 0.40307f
C5918 a_5396_8177.t35 AVSS 0.095293f
C5919 a_5396_8177.t5 AVSS 0.095293f
C5920 a_5396_8177.n71 AVSS 0.411692f
C5921 a_5396_8177.t67 AVSS 0.403593f
C5922 a_5396_8177.t20 AVSS 0.403593f
C5923 a_5396_8177.n72 AVSS 0.265627f
C5924 a_5396_8177.n73 AVSS 3.88765f
C5925 a_5396_8177.n74 AVSS 6.4282f
C5926 a_5396_8177.t15 AVSS 0.538544f
C5927 a_5396_8177.t8 AVSS 0.095293f
C5928 a_5396_8177.t46 AVSS 0.095293f
C5929 a_5396_8177.n75 AVSS 0.411692f
C5930 a_5396_8177.t42 AVSS 0.403593f
C5931 a_5396_8177.t78 AVSS 0.40307f
C5932 a_5396_8177.t16 AVSS 0.095293f
C5933 a_5396_8177.t10 AVSS 0.095293f
C5934 a_5396_8177.n76 AVSS 0.411692f
C5935 a_5396_8177.t37 AVSS 0.403593f
C5936 a_5396_8177.t62 AVSS 0.403593f
C5937 a_5396_8177.t57 AVSS 0.095293f
C5938 a_5396_8177.t82 AVSS 0.095293f
C5939 a_5396_8177.n77 AVSS 0.411692f
C5940 a_5396_8177.t79 AVSS 0.403593f
C5941 a_5396_8177.t7 AVSS 0.40307f
C5942 a_5396_8177.t36 AVSS 0.095293f
C5943 a_5396_8177.t30 AVSS 0.095293f
C5944 a_5396_8177.n78 AVSS 0.411692f
C5945 a_5396_8177.t77 AVSS 0.539266f
C5946 a_5396_8177.n79 AVSS 3.81741f
C5947 a_5396_8177.t88 AVSS 0.095293f
C5948 a_5396_8177.t170 AVSS 0.095293f
C5949 a_5396_8177.n80 AVSS 0.523527f
C5950 a_5396_8177.t121 AVSS 0.095293f
C5951 a_5396_8177.t118 AVSS 0.095293f
C5952 a_5396_8177.n81 AVSS 0.349599f
C5953 a_5396_8177.n82 AVSS 1.7194f
C5954 a_5396_8177.t150 AVSS 0.095293f
C5955 a_5396_8177.t90 AVSS 0.095293f
C5956 a_5396_8177.n83 AVSS 0.349599f
C5957 a_5396_8177.n84 AVSS 1.21944f
C5958 a_5396_8177.t172 AVSS 0.095293f
C5959 a_5396_8177.t110 AVSS 0.095293f
C5960 a_5396_8177.n85 AVSS 0.349599f
C5961 a_5396_8177.n86 AVSS 0.489773f
C5962 a_5396_8177.n87 AVSS 4.03456f
C5963 a_5396_8177.t175 AVSS 0.095293f
C5964 a_5396_8177.t113 AVSS 0.095293f
C5965 a_5396_8177.n88 AVSS 0.522186f
C5966 a_5396_8177.t148 AVSS 0.095293f
C5967 a_5396_8177.t119 AVSS 0.095293f
C5968 a_5396_8177.n89 AVSS 0.348584f
C5969 a_5396_8177.t116 AVSS 0.095293f
C5970 a_5396_8177.t144 AVSS 0.095293f
C5971 a_5396_8177.n90 AVSS 0.348584f
C5972 a_5396_8177.t94 AVSS 0.095293f
C5973 a_5396_8177.t127 AVSS 0.095293f
C5974 a_5396_8177.n91 AVSS 0.348584f
C5975 a_5396_8177.t137 AVSS 0.095293f
C5976 a_5396_8177.t100 AVSS 0.095293f
C5977 a_5396_8177.n92 AVSS 0.348584f
C5978 a_5396_8177.t115 AVSS 0.095293f
C5979 a_5396_8177.t164 AVSS 0.095293f
C5980 a_5396_8177.n93 AVSS 0.348584f
C5981 a_5396_8177.t160 AVSS 0.095293f
C5982 a_5396_8177.t108 AVSS 0.095293f
C5983 a_5396_8177.n94 AVSS 0.348584f
C5984 a_5396_8177.t158 AVSS 0.095293f
C5985 a_5396_8177.t171 AVSS 0.095293f
C5986 a_5396_8177.n95 AVSS 0.348584f
C5987 a_5396_8177.t106 AVSS 0.095293f
C5988 a_5396_8177.t162 AVSS 0.095293f
C5989 a_5396_8177.n96 AVSS 0.262891f
C5990 a_5396_8177.t105 AVSS 0.095293f
C5991 a_5396_8177.t161 AVSS 0.095293f
C5992 a_5396_8177.n97 AVSS 0.240067f
C5993 a_5396_8177.n98 AVSS 1.47694f
C5994 a_5396_8177.t143 AVSS 0.268949f
C5995 a_5396_8177.t142 AVSS 0.249568f
C5996 a_5396_8177.n99 AVSS 0.855341f
C5997 a_5396_8177.n100 AVSS 1.6948f
C5998 a_5396_8177.t167 AVSS 0.095293f
C5999 a_5396_8177.t147 AVSS 0.095293f
C6000 a_5396_8177.n101 AVSS 0.522186f
C6001 a_5396_8177.t131 AVSS 0.095293f
C6002 a_5396_8177.t112 AVSS 0.095293f
C6003 a_5396_8177.n102 AVSS 0.348584f
C6004 a_5396_8177.t135 AVSS 0.095293f
C6005 a_5396_8177.t104 AVSS 0.095293f
C6006 a_5396_8177.n103 AVSS 0.348584f
C6007 a_5396_8177.t163 AVSS 0.095293f
C6008 a_5396_8177.t139 AVSS 0.095293f
C6009 a_5396_8177.n104 AVSS 0.348584f
C6010 a_5396_8177.t91 AVSS 0.095293f
C6011 a_5396_8177.t157 AVSS 0.095293f
C6012 a_5396_8177.n105 AVSS 0.348584f
C6013 a_5396_8177.t122 AVSS 0.095293f
C6014 a_5396_8177.t101 AVSS 0.095293f
C6015 a_5396_8177.n106 AVSS 0.348584f
C6016 a_5396_8177.t140 AVSS 0.095293f
C6017 a_5396_8177.t114 AVSS 0.095293f
C6018 a_5396_8177.n107 AVSS 0.348584f
C6019 a_5396_8177.t96 AVSS 0.095293f
C6020 a_5396_8177.t126 AVSS 0.095293f
C6021 a_5396_8177.n108 AVSS 0.348584f
C6022 a_5396_8177.n109 AVSS 1.64011f
C6023 a_5396_8177.n110 AVSS 5.54716f
C6024 a_5396_8177.n111 AVSS 1.80856f
C6025 a_5396_8177.t95 AVSS 0.095293f
C6026 a_5396_8177.t154 AVSS 0.095293f
C6027 a_5396_8177.n112 AVSS 0.262891f
C6028 a_5396_8177.t93 AVSS 0.095293f
C6029 a_5396_8177.t153 AVSS 0.095293f
C6030 a_5396_8177.n113 AVSS 0.240067f
C6031 a_5396_8177.n114 AVSS 0.662164f
C6032 a_5396_8177.n115 AVSS 1.57141f
C6033 a_5396_8177.t134 AVSS 0.268949f
C6034 a_5396_8177.t133 AVSS 0.249568f
C6035 a_5396_8177.n116 AVSS 0.855341f
C6036 a_5396_8177.n117 AVSS 1.02367f
C6037 a_5396_8177.n118 AVSS 6.10479f
C6038 a_5396_8177.t155 AVSS 0.095293f
C6039 a_5396_8177.t138 AVSS 0.095293f
C6040 a_5396_8177.n119 AVSS 0.523527f
C6041 a_5396_8177.t117 AVSS 0.095293f
C6042 a_5396_8177.t97 AVSS 0.095293f
C6043 a_5396_8177.n120 AVSS 0.349599f
C6044 a_5396_8177.n121 AVSS 1.7194f
C6045 a_5396_8177.t120 AVSS 0.095293f
C6046 a_5396_8177.t92 AVSS 0.095293f
C6047 a_5396_8177.n122 AVSS 0.349599f
C6048 a_5396_8177.n123 AVSS 1.21944f
C6049 a_5396_8177.t151 AVSS 0.095293f
C6050 a_5396_8177.t123 AVSS 0.095293f
C6051 a_5396_8177.n124 AVSS 0.349599f
C6052 a_5396_8177.n125 AVSS 0.489773f
C6053 a_5396_8177.n126 AVSS 0.794685f
C6054 a_5396_8177.t159 AVSS 0.095293f
C6055 a_5396_8177.t141 AVSS 0.095293f
C6056 a_5396_8177.n127 AVSS 0.349599f
C6057 a_5396_8177.n128 AVSS 1.18797f
C6058 a_5396_8177.t107 AVSS 0.095293f
C6059 a_5396_8177.t89 AVSS 0.095293f
C6060 a_5396_8177.n129 AVSS 0.349599f
C6061 a_5396_8177.n130 AVSS 1.21941f
C6062 a_5396_8177.t130 AVSS 0.095293f
C6063 a_5396_8177.t98 AVSS 0.095293f
C6064 a_5396_8177.n131 AVSS 0.349599f
C6065 a_5396_8177.n132 AVSS 1.21944f
C6066 a_5396_8177.t165 AVSS 0.095293f
C6067 a_5396_8177.t111 AVSS 0.095293f
C6068 a_5396_8177.n133 AVSS 0.349599f
C6069 a_5396_8177.n134 AVSS 0.749824f
C6070 a_5396_8177.n135 AVSS 4.0754f
C6071 a_5396_8177.n136 AVSS 3.92753f
C6072 a_5396_8177.n137 AVSS 0.794608f
C6073 a_5396_8177.n138 AVSS 3.88513f
C6074 a_5396_8177.t145 AVSS 0.095293f
C6075 a_5396_8177.t173 AVSS 0.095293f
C6076 a_5396_8177.n139 AVSS 0.262891f
C6077 a_5396_8177.t146 AVSS 0.095293f
C6078 a_5396_8177.t174 AVSS 0.095293f
C6079 a_5396_8177.n140 AVSS 0.240067f
C6080 a_5396_8177.n141 AVSS 1.47694f
C6081 a_5396_8177.t166 AVSS 0.268949f
C6082 a_5396_8177.t168 AVSS 0.249568f
C6083 a_5396_8177.n142 AVSS 0.855341f
C6084 a_5396_8177.n143 AVSS 1.6948f
C6085 a_5396_8177.t124 AVSS 0.268949f
C6086 a_5396_8177.t125 AVSS 0.249568f
C6087 a_5396_8177.n144 AVSS 0.855341f
C6088 a_5396_8177.n145 AVSS 1.02367f
C6089 a_5396_8177.t99 AVSS 0.095293f
C6090 a_5396_8177.t128 AVSS 0.095293f
C6091 a_5396_8177.n146 AVSS 0.262891f
C6092 a_5396_8177.t102 AVSS 0.095293f
C6093 a_5396_8177.t129 AVSS 0.095293f
C6094 a_5396_8177.n147 AVSS 0.240067f
C6095 a_5396_8177.n148 AVSS 0.662164f
C6096 a_5396_8177.n149 AVSS 1.57141f
C6097 a_5396_8177.n150 AVSS 1.80856f
C6098 a_5396_8177.n151 AVSS 3.37808f
C6099 a_5396_8177.n152 AVSS 4.68889f
C6100 a_5396_8177.n153 AVSS 0.794685f
C6101 a_5396_8177.t136 AVSS 0.095293f
C6102 a_5396_8177.t132 AVSS 0.095293f
C6103 a_5396_8177.n154 AVSS 0.349599f
C6104 a_5396_8177.n155 AVSS 1.18797f
C6105 a_5396_8177.t156 AVSS 0.095293f
C6106 a_5396_8177.t152 AVSS 0.095293f
C6107 a_5396_8177.n156 AVSS 0.349599f
C6108 a_5396_8177.n157 AVSS 1.21941f
C6109 a_5396_8177.t169 AVSS 0.095293f
C6110 a_5396_8177.t109 AVSS 0.095293f
C6111 a_5396_8177.n158 AVSS 0.349599f
C6112 a_5396_8177.n159 AVSS 1.21944f
C6113 a_5396_8177.t103 AVSS 0.095293f
C6114 a_5396_8177.t149 AVSS 0.095293f
C6115 a_5396_8177.n160 AVSS 0.349599f
C6116 a_5396_8177.n161 AVSS 0.749824f
C6117 a_5396_8177.n162 AVSS 5.24322f
C6118 a_5396_8177.n163 AVSS 6.28145f
C6119 a_5396_8177.n164 AVSS 4.10788f
C6120 a_5396_8177.n165 AVSS 0.265627f
C6121 a_5396_8177.n166 AVSS 0.265627f
C6122 a_5396_8177.n167 AVSS 4.55647f
C6123 a_5396_8177.t60 AVSS 0.234869f
C6124 a_5396_8177.t3 AVSS 0.28657f
C6125 a_5396_8177.n168 AVSS 1.53577f
C6126 a_5396_8177.t31 AVSS 0.095293f
C6127 a_5396_8177.t13 AVSS 0.095293f
C6128 a_5396_8177.n169 AVSS 0.22302f
C6129 a_5396_8177.t27 AVSS 0.095293f
C6130 a_5396_8177.t23 AVSS 0.095293f
C6131 a_5396_8177.n170 AVSS 0.283728f
C6132 a_5396_8177.n171 AVSS 0.645783f
C6133 a_5396_8177.n172 AVSS 1.41165f
C6134 a_5396_8177.t19 AVSS 0.095293f
C6135 a_5396_8177.t86 AVSS 0.095293f
C6136 a_5396_8177.n173 AVSS 0.22302f
C6137 a_5396_8177.t70 AVSS 0.095293f
C6138 a_5396_8177.t65 AVSS 0.095293f
C6139 a_5396_8177.n174 AVSS 0.283728f
C6140 a_5396_8177.n175 AVSS 0.645783f
C6141 a_5396_8177.n176 AVSS 1.12242f
C6142 a_5396_8177.t48 AVSS 0.234869f
C6143 a_5396_8177.t43 AVSS 0.28657f
C6144 a_5396_8177.n177 AVSS 0.839828f
C6145 a_5396_8177.n178 AVSS 1.71657f
C6146 a_5396_8177.n179 AVSS 1.80896f
C6147 a_5396_8177.n180 AVSS 3.91535f
C6148 a_5396_8177.n181 AVSS 3.49477f
C6149 a_5396_8177.n182 AVSS 0.265638f
C6150 a_5396_8177.t59 AVSS 0.095293f
C6151 a_5396_8177.t34 AVSS 0.095293f
C6152 a_5396_8177.n183 AVSS 0.41253f
C6153 a_5396_8177.n184 AVSS 0.619074f
C6154 a_5396_8177.t4 AVSS 0.404302f
C6155 a_5396_8177.n185 AVSS 1.16606f
C6156 a_5396_8177.t45 AVSS 0.400953f
C6157 a_5396_8177.n186 AVSS 1.15658f
C6158 a_5396_8177.t26 AVSS 0.095293f
C6159 a_5396_8177.t75 AVSS 0.095293f
C6160 a_5396_8177.n187 AVSS 0.41253f
C6161 a_5396_8177.n188 AVSS 0.78412f
C6162 a_5396_8177.t56 AVSS 0.404415f
C6163 a_5396_8177.n189 AVSS 1.14932f
C6164 a_5396_8177.t9 AVSS 0.400953f
C6165 a_5396_8177.n190 AVSS 1.04137f
C6166 a_5396_8177.t80 AVSS 0.541038f
C6167 a_5396_8177.t71 AVSS 0.095293f
C6168 a_5396_8177.t49 AVSS 0.095293f
C6169 a_5396_8177.n191 AVSS 0.41253f
C6170 a_5396_8177.n192 AVSS 1.21102f
C6171 a_5396_8177.n193 AVSS 0.265638f
C6172 a_5396_8177.n194 AVSS 3.49477f
C6173 a_5396_8177.n195 AVSS 3.88765f
C6174 a_5396_8177.n196 AVSS 0.265627f
C6175 a_5396_8177.n197 AVSS 0.411692f
C6176 a_5396_8177.t87 AVSS 0.095293f
C6177 a_5396_n6451.n0 AVSS 0.519739f
C6178 a_5396_n6451.n1 AVSS 0.967963f
C6179 a_5396_n6451.n2 AVSS 1.05403f
C6180 a_5396_n6451.n3 AVSS 0.967963f
C6181 a_5396_n6451.n4 AVSS 1.05403f
C6182 a_5396_n6451.n5 AVSS 0.988808f
C6183 a_5396_n6451.n6 AVSS 1.50233f
C6184 a_5396_n6451.n7 AVSS 0.772166f
C6185 a_5396_n6451.n8 AVSS 1.04659f
C6186 a_5396_n6451.n9 AVSS 0.393209f
C6187 a_5396_n6451.n10 AVSS 1.04659f
C6188 a_5396_n6451.n11 AVSS 0.772166f
C6189 a_5396_n6451.n12 AVSS 0.390068f
C6190 a_5396_n6451.n13 AVSS 1.35517f
C6191 a_5396_n6451.n14 AVSS 0.988167f
C6192 a_5396_n6451.n15 AVSS 0.388938f
C6193 a_5396_n6451.n16 AVSS 1.05523f
C6194 a_5396_n6451.n17 AVSS 0.769779f
C6195 a_5396_n6451.n18 AVSS 0.56328f
C6196 a_5396_n6451.n19 AVSS 0.294838f
C6197 a_5396_n6451.n20 AVSS 0.609323f
C6198 a_5396_n6451.n21 AVSS 0.72635f
C6199 a_5396_n6451.n22 AVSS 0.988167f
C6200 a_5396_n6451.n23 AVSS 1.35517f
C6201 a_5396_n6451.n24 AVSS 0.56328f
C6202 a_5396_n6451.n25 AVSS 0.769779f
C6203 a_5396_n6451.n26 AVSS 1.05523f
C6204 a_5396_n6451.n27 AVSS 1.45171f
C6205 a_5396_n6451.n28 AVSS 0.963935f
C6206 a_5396_n6451.n29 AVSS 1.0503f
C6207 a_5396_n6451.n30 AVSS 0.963935f
C6208 a_5396_n6451.n31 AVSS 1.0503f
C6209 a_5396_n6451.n32 AVSS 0.716301f
C6210 a_5396_n6451.n33 AVSS 0.988808f
C6211 a_5396_n6451.n34 AVSS 1.34487f
C6212 a_5396_n6451.n35 AVSS 0.39289f
C6213 a_5396_n6451.n36 AVSS 1.34487f
C6214 a_5396_n6451.n37 AVSS 0.388938f
C6215 a_5396_n6451.n38 AVSS 0.74452f
C6216 a_5396_n6451.n39 AVSS 0.388938f
C6217 a_5396_n6451.n40 AVSS 0.609323f
C6218 a_5396_n6451.n41 AVSS 0.74452f
C6219 a_5396_n6451.n42 AVSS 0.294838f
C6220 a_5396_n6451.n43 AVSS 0.599334f
C6221 a_5396_n6451.n44 AVSS 0.569992f
C6222 a_5396_n6451.n45 AVSS 0.750301f
C6223 a_5396_n6451.n46 AVSS 0.599334f
C6224 a_5396_n6451.n47 AVSS 0.716301f
C6225 a_5396_n6451.n48 AVSS 0.393209f
C6226 a_5396_n6451.n49 AVSS 0.296095f
C6227 a_5396_n6451.n50 AVSS 0.393209f
C6228 a_5396_n6451.n51 AVSS 0.750301f
C6229 a_5396_n6451.n52 AVSS 0.296095f
C6230 a_5396_n6451.n53 AVSS 0.612855f
C6231 a_5396_n6451.n54 AVSS 0.854088f
C6232 a_5396_n6451.n55 AVSS 2.60496f
C6233 a_5396_n6451.n56 AVSS 0.946222f
C6234 a_5396_n6451.n57 AVSS 0.667759f
C6235 a_5396_n6451.n58 AVSS 1.05756f
C6236 a_5396_n6451.n59 AVSS 2.60496f
C6237 a_5396_n6451.n60 AVSS 0.9706f
C6238 a_5396_n6451.n61 AVSS 0.9706f
C6239 a_5396_n6451.n62 AVSS 0.946222f
C6240 a_5396_n6451.n63 AVSS 2.60496f
C6241 a_5396_n6451.n64 AVSS 0.854088f
C6242 a_5396_n6451.n65 AVSS 1.1094f
C6243 a_5396_n6451.n66 AVSS 1.85373f
C6244 a_5396_n6451.n67 AVSS 0.64731f
C6245 a_5396_n6451.n68 AVSS 2.60496f
C6246 a_5396_n6451.n69 AVSS 1.05756f
C6247 a_5396_n6451.n70 AVSS 1.35705f
C6248 a_5396_n6451.n71 AVSS 1.3878f
C6249 a_5396_n6451.n72 AVSS 2.654f
C6250 a_5396_n6451.n73 AVSS 1.04821f
C6251 a_5396_n6451.n74 AVSS 0.879243f
C6252 a_5396_n6451.n75 AVSS 2.64918f
C6253 a_5396_n6451.n76 AVSS 0.923787f
C6254 a_5396_n6451.n77 AVSS 1.1119f
C6255 a_5396_n6451.n78 AVSS 1.93453f
C6256 a_5396_n6451.n79 AVSS 0.686793f
C6257 a_5396_n6451.n80 AVSS 0.976242f
C6258 a_5396_n6451.n81 AVSS 0.623461f
C6259 a_5396_n6451.n82 AVSS 1.04818f
C6260 a_5396_n6451.n83 AVSS 0.879251f
C6261 a_5396_n6451.n84 AVSS 0.923788f
C6262 a_5396_n6451.n85 AVSS 2.64918f
C6263 a_5396_n6451.n86 AVSS 2.654f
C6264 a_5396_n6451.n87 AVSS 0.976215f
C6265 a_5396_n6451.n88 AVSS 0.72635f
C6266 a_5396_n6451.n89 AVSS 1.85373f
C6267 a_5396_n6451.n90 AVSS 0.64817f
C6268 a_5396_n6451.n91 AVSS 1.85373f
C6269 a_5396_n6451.n92 AVSS 0.64731f
C6270 a_5396_n6451.n93 AVSS 1.85373f
C6271 a_5396_n6451.n94 AVSS 0.64817f
C6272 a_5396_n6451.n95 AVSS 1.3635f
C6273 a_5396_n6451.n96 AVSS 2.51808f
C6274 a_5396_n6451.n97 AVSS 2.51808f
C6275 a_5396_n6451.n98 AVSS 1.3635f
C6276 a_5396_n6451.n99 AVSS 1.93453f
C6277 a_5396_n6451.n100 AVSS 0.686801f
C6278 a_5396_n6451.n101 AVSS 1.93453f
C6279 a_5396_n6451.n102 AVSS 0.638702f
C6280 a_5396_n6451.n103 AVSS 1.93453f
C6281 a_5396_n6451.n104 AVSS 0.638684f
C6282 a_5396_n6451.n105 AVSS 1.38647f
C6283 a_5396_n6451.n106 AVSS 2.54499f
C6284 a_5396_n6451.n107 AVSS 2.54499f
C6285 a_5396_n6451.n108 AVSS 1.38647f
C6286 a_5396_n6451.n109 AVSS 1.1094f
C6287 a_5396_n6451.n110 AVSS 2.51711f
C6288 a_5396_n6451.n111 AVSS 0.667759f
C6289 a_5396_n6451.n112 AVSS 2.51711f
C6290 a_5396_n6451.n113 AVSS 0.654202f
C6291 a_5396_n6451.n114 AVSS 1.1119f
C6292 a_5396_n6451.n115 AVSS 2.53269f
C6293 a_5396_n6451.n116 AVSS 2.53269f
C6294 a_5396_n6451.n117 AVSS 0.612855f
C6295 a_5396_n6451.t167 AVSS 0.532372f
C6296 a_5396_n6451.t242 AVSS 0.532372f
C6297 a_5396_n6451.n118 AVSS 0.812058f
C6298 a_5396_n6451.n119 AVSS 0.634079f
C6299 a_5396_n6451.n120 AVSS 0.695469f
C6300 a_5396_n6451.n121 AVSS 0.557171f
C6301 a_5396_n6451.n122 AVSS 0.70564f
C6302 a_5396_n6451.n123 AVSS 0.705639f
C6303 a_5396_n6451.n124 AVSS 0.456781f
C6304 a_5396_n6451.n125 AVSS 0.634079f
C6305 a_5396_n6451.n126 AVSS 0.695469f
C6306 a_5396_n6451.n127 AVSS 0.910589f
C6307 a_5396_n6451.n128 AVSS 0.812058f
C6308 a_5396_n6451.n129 AVSS 0.634079f
C6309 a_5396_n6451.n130 AVSS 0.695469f
C6310 a_5396_n6451.n131 AVSS 0.557171f
C6311 a_5396_n6451.n132 AVSS 0.70564f
C6312 a_5396_n6451.n133 AVSS 0.705639f
C6313 a_5396_n6451.n134 AVSS 0.456781f
C6314 a_5396_n6451.n135 AVSS 0.634079f
C6315 a_5396_n6451.n136 AVSS 0.695469f
C6316 a_5396_n6451.n137 AVSS 0.910589f
C6317 a_5396_n6451.n138 AVSS 1.16738f
C6318 a_5396_n6451.t17 AVSS 0.825042f
C6319 a_5396_n6451.t8 AVSS 0.24494f
C6320 a_5396_n6451.n139 AVSS 0.905519f
C6321 a_5396_n6451.n140 AVSS 2.39697f
C6322 a_5396_n6451.n141 AVSS 2.14352f
C6323 a_5396_n6451.n142 AVSS 2.35461f
C6324 a_5396_n6451.t52 AVSS 1.08015f
C6325 a_5396_n6451.n143 AVSS 2.37139f
C6326 a_5396_n6451.t16 AVSS 3.04535f
C6327 a_5396_n6451.n144 AVSS 3.42133f
C6328 a_5396_n6451.t226 AVSS 0.481683f
C6329 a_5396_n6451.t216 AVSS 0.530966f
C6330 a_5396_n6451.t147 AVSS 0.481683f
C6331 a_5396_n6451.t155 AVSS 0.481683f
C6332 a_5396_n6451.t237 AVSS 0.481683f
C6333 a_5396_n6451.n145 AVSS 0.390068f
C6334 a_5396_n6451.t185 AVSS 0.481683f
C6335 a_5396_n6451.n146 AVSS 0.320727f
C6336 a_5396_n6451.t193 AVSS 0.481683f
C6337 a_5396_n6451.t223 AVSS 0.481683f
C6338 a_5396_n6451.t168 AVSS 0.481683f
C6339 a_5396_n6451.t125 AVSS 0.481683f
C6340 a_5396_n6451.t77 AVSS 0.481683f
C6341 a_5396_n6451.t85 AVSS 0.481683f
C6342 a_5396_n6451.t202 AVSS 0.481683f
C6343 a_5396_n6451.t172 AVSS 0.481683f
C6344 a_5396_n6451.t113 AVSS 0.481683f
C6345 a_5396_n6451.t162 AVSS 0.481683f
C6346 a_5396_n6451.t123 AVSS 0.481683f
C6347 a_5396_n6451.t83 AVSS 0.481683f
C6348 a_5396_n6451.t221 AVSS 0.530966f
C6349 a_5396_n6451.t105 AVSS 0.481683f
C6350 a_5396_n6451.t145 AVSS 0.481683f
C6351 a_5396_n6451.t184 AVSS 0.481683f
C6352 a_5396_n6451.t192 AVSS 0.481683f
C6353 a_5396_n6451.n147 AVSS 0.39289f
C6354 a_5396_n6451.t76 AVSS 0.481683f
C6355 a_5396_n6451.n148 AVSS 0.320727f
C6356 a_5396_n6451.t114 AVSS 0.481683f
C6357 a_5396_n6451.t195 AVSS 0.481683f
C6358 a_5396_n6451.t73 AVSS 0.481683f
C6359 a_5396_n6451.t89 AVSS 0.481683f
C6360 a_5396_n6451.t161 AVSS 0.481683f
C6361 a_5396_n6451.t199 AVSS 0.481683f
C6362 a_5396_n6451.t116 AVSS 0.481683f
C6363 a_5396_n6451.t174 AVSS 0.481683f
C6364 a_5396_n6451.t217 AVSS 0.481683f
C6365 a_5396_n6451.t156 AVSS 0.532447f
C6366 a_5396_n6451.t139 AVSS 0.481683f
C6367 a_5396_n6451.n149 AVSS 0.393209f
C6368 a_5396_n6451.t98 AVSS 0.481683f
C6369 a_5396_n6451.n150 AVSS 0.320727f
C6370 a_5396_n6451.t220 AVSS 0.481683f
C6371 a_5396_n6451.t228 AVSS 0.481683f
C6372 a_5396_n6451.t131 AVSS 0.481683f
C6373 a_5396_n6451.t136 AVSS 0.481683f
C6374 a_5396_n6451.n151 AVSS 5.14918f
C6375 a_5396_n6451.n152 AVSS 0.519739f
C6376 a_5396_n6451.t182 AVSS 0.481683f
C6377 a_5396_n6451.n153 AVSS 0.390068f
C6378 a_5396_n6451.t241 AVSS 0.481683f
C6379 a_5396_n6451.n154 AVSS 0.320727f
C6380 a_5396_n6451.t104 AVSS 0.481683f
C6381 a_5396_n6451.t229 AVSS 0.481683f
C6382 a_5396_n6451.t109 AVSS 0.481683f
C6383 a_5396_n6451.t67 AVSS 0.481683f
C6384 a_5396_n6451.t138 AVSS 0.481683f
C6385 a_5396_n6451.t176 AVSS 0.481683f
C6386 a_5396_n6451.t210 AVSS 0.481683f
C6387 a_5396_n6451.n155 AVSS 0.390068f
C6388 a_5396_n6451.t93 AVSS 0.481683f
C6389 a_5396_n6451.n156 AVSS 0.320727f
C6390 a_5396_n6451.t129 AVSS 0.481683f
C6391 a_5396_n6451.t134 AVSS 0.533378f
C6392 a_5396_n6451.t191 AVSS 0.481683f
C6393 a_5396_n6451.t151 AVSS 0.481683f
C6394 a_5396_n6451.t95 AVSS 0.481683f
C6395 a_5396_n6451.n157 AVSS 5.14918f
C6396 a_5396_n6451.t238 AVSS 0.481683f
C6397 a_5396_n6451.n158 AVSS 0.519371f
C6398 a_5396_n6451.t111 AVSS 0.481683f
C6399 a_5396_n6451.t208 AVSS 0.481683f
C6400 a_5396_n6451.t74 AVSS 0.481683f
C6401 a_5396_n6451.t120 AVSS 0.481683f
C6402 a_5396_n6451.n159 AVSS 0.39289f
C6403 a_5396_n6451.t178 AVSS 0.481683f
C6404 a_5396_n6451.n160 AVSS 0.320727f
C6405 a_5396_n6451.t219 AVSS 0.481683f
C6406 a_5396_n6451.t121 AVSS 0.481683f
C6407 a_5396_n6451.t173 AVSS 0.481683f
C6408 a_5396_n6451.t233 AVSS 0.481683f
C6409 a_5396_n6451.t150 AVSS 0.481683f
C6410 a_5396_n6451.t188 AVSS 0.481683f
C6411 a_5396_n6451.t92 AVSS 0.481683f
C6412 a_5396_n6451.t128 AVSS 0.481683f
C6413 a_5396_n6451.t144 AVSS 0.481683f
C6414 a_5396_n6451.n161 AVSS 0.39289f
C6415 a_5396_n6451.t204 AVSS 0.481683f
C6416 a_5396_n6451.n162 AVSS 0.320727f
C6417 a_5396_n6451.t68 AVSS 0.481683f
C6418 a_5396_n6451.t101 AVSS 0.481683f
C6419 a_5396_n6451.t141 AVSS 0.481683f
C6420 a_5396_n6451.t84 AVSS 0.532447f
C6421 a_5396_n6451.t224 AVSS 0.481683f
C6422 a_5396_n6451.n163 AVSS 3.42133f
C6423 a_5396_n6451.n164 AVSS 3.65785f
C6424 a_5396_n6451.t227 AVSS 0.481683f
C6425 a_5396_n6451.t171 AVSS 0.481683f
C6426 a_5396_n6451.t180 AVSS 0.481683f
C6427 a_5396_n6451.t88 AVSS 0.533378f
C6428 a_5396_n6451.t112 AVSS 0.481683f
C6429 a_5396_n6451.n165 AVSS 0.388938f
C6430 a_5396_n6451.t102 AVSS 0.481683f
C6431 a_5396_n6451.n166 AVSS 0.320727f
C6432 a_5396_n6451.t153 AVSS 0.481683f
C6433 a_5396_n6451.t115 AVSS 0.481683f
C6434 a_5396_n6451.t213 AVSS 0.481683f
C6435 a_5396_n6451.t86 AVSS 0.481683f
C6436 a_5396_n6451.n167 AVSS 3.65785f
C6437 a_5396_n6451.n168 AVSS 2.83294f
C6438 a_5396_n6451.n169 AVSS 3.42133f
C6439 a_5396_n6451.t169 AVSS 0.481683f
C6440 a_5396_n6451.t236 AVSS 0.481683f
C6441 a_5396_n6451.t110 AVSS 0.481683f
C6442 a_5396_n6451.t206 AVSS 0.481683f
C6443 a_5396_n6451.t194 AVSS 0.481683f
C6444 a_5396_n6451.t154 AVSS 0.481683f
C6445 a_5396_n6451.t148 AVSS 0.481683f
C6446 a_5396_n6451.t108 AVSS 0.481683f
C6447 a_5396_n6451.t70 AVSS 0.481683f
C6448 a_5396_n6451.t187 AVSS 0.481683f
C6449 a_5396_n6451.t215 AVSS 0.481683f
C6450 a_5396_n6451.t78 AVSS 0.481683f
C6451 a_5396_n6451.t197 AVSS 0.481683f
C6452 a_5396_n6451.t80 AVSS 0.481683f
C6453 a_5396_n6451.t135 AVSS 0.481683f
C6454 a_5396_n6451.t165 AVSS 0.481683f
C6455 a_5396_n6451.t203 AVSS 0.481683f
C6456 a_5396_n6451.t146 AVSS 0.481683f
C6457 a_5396_n6451.t214 AVSS 0.481683f
C6458 a_5396_n6451.t149 AVSS 0.481683f
C6459 a_5396_n6451.t177 AVSS 0.481683f
C6460 a_5396_n6451.t198 AVSS 0.481683f
C6461 a_5396_n6451.t160 AVSS 0.481683f
C6462 a_5396_n6451.t82 AVSS 0.481683f
C6463 a_5396_n6451.t119 AVSS 0.481683f
C6464 a_5396_n6451.t235 AVSS 0.481683f
C6465 a_5396_n6451.t97 AVSS 0.481683f
C6466 a_5396_n6451.t90 AVSS 0.481683f
C6467 a_5396_n6451.t240 AVSS 0.481683f
C6468 a_5396_n6451.t103 AVSS 0.481683f
C6469 a_5396_n6451.t175 AVSS 0.481683f
C6470 a_5396_n6451.t218 AVSS 0.481683f
C6471 a_5396_n6451.t87 AVSS 0.481683f
C6472 a_5396_n6451.t124 AVSS 0.481683f
C6473 a_5396_n6451.t133 AVSS 0.481683f
C6474 a_5396_n6451.t190 AVSS 0.481683f
C6475 a_5396_n6451.t231 AVSS 0.481683f
C6476 a_5396_n6451.t170 AVSS 0.481683f
C6477 a_5396_n6451.n170 AVSS 5.34741f
C6478 a_5396_n6451.t205 AVSS 0.481683f
C6479 a_5396_n6451.t239 AVSS 0.481683f
C6480 a_5396_n6451.t99 AVSS 0.481683f
C6481 a_5396_n6451.t122 AVSS 0.481683f
C6482 a_5396_n6451.t179 AVSS 0.481683f
C6483 a_5396_n6451.t222 AVSS 0.481683f
C6484 a_5396_n6451.t159 AVSS 0.481683f
C6485 a_5396_n6451.t181 AVSS 0.481683f
C6486 a_5396_n6451.t94 AVSS 0.481683f
C6487 a_5396_n6451.t232 AVSS 0.481683f
C6488 a_5396_n6451.t142 AVSS 0.481683f
C6489 a_5396_n6451.n171 AVSS 5.34741f
C6490 a_5396_n6451.t107 AVSS 0.481683f
C6491 a_5396_n6451.t183 AVSS 0.481683f
C6492 a_5396_n6451.t225 AVSS 0.481683f
C6493 a_5396_n6451.t91 AVSS 0.481683f
C6494 a_5396_n6451.t126 AVSS 0.481683f
C6495 a_5396_n6451.t163 AVSS 0.481683f
C6496 a_5396_n6451.t201 AVSS 0.481683f
C6497 a_5396_n6451.t81 AVSS 0.481683f
C6498 a_5396_n6451.t137 AVSS 0.481683f
C6499 a_5396_n6451.t189 AVSS 0.481683f
C6500 a_5396_n6451.t75 AVSS 0.481683f
C6501 a_5396_n6451.t186 AVSS 0.481683f
C6502 a_5396_n6451.t230 AVSS 0.481683f
C6503 a_5396_n6451.t234 AVSS 0.481683f
C6504 a_5396_n6451.t117 AVSS 0.481683f
C6505 a_5396_n6451.t157 AVSS 0.481683f
C6506 a_5396_n6451.t96 AVSS 0.481683f
C6507 a_5396_n6451.t130 AVSS 0.481683f
C6508 a_5396_n6451.t143 AVSS 0.481683f
C6509 a_5396_n6451.t106 AVSS 0.481683f
C6510 a_5396_n6451.t207 AVSS 0.481683f
C6511 a_5396_n6451.t166 AVSS 0.481683f
C6512 a_5396_n6451.n172 AVSS 3.42133f
C6513 a_5396_n6451.n173 AVSS 3.88032f
C6514 a_5396_n6451.t79 AVSS 0.481683f
C6515 a_5396_n6451.t140 AVSS 0.481683f
C6516 a_5396_n6451.t132 AVSS 0.481683f
C6517 a_5396_n6451.t209 AVSS 0.481683f
C6518 a_5396_n6451.t196 AVSS 0.481683f
C6519 a_5396_n6451.t200 AVSS 0.481683f
C6520 a_5396_n6451.t212 AVSS 0.481683f
C6521 a_5396_n6451.t71 AVSS 0.481683f
C6522 a_5396_n6451.t152 AVSS 0.481683f
C6523 a_5396_n6451.t100 AVSS 0.481683f
C6524 a_5396_n6451.t69 AVSS 0.481683f
C6525 a_5396_n6451.t118 AVSS 0.481683f
C6526 a_5396_n6451.t127 AVSS 0.481683f
C6527 a_5396_n6451.t158 AVSS 0.481683f
C6528 a_5396_n6451.t164 AVSS 0.481683f
C6529 a_5396_n6451.t72 AVSS 0.481683f
C6530 a_5396_n6451.t211 AVSS 0.481683f
C6531 a_5396_n6451.n174 AVSS 3.48859f
C6532 a_5396_n6451.n175 AVSS 3.51576f
C6533 a_5396_n6451.n176 AVSS 2.65516f
C6534 a_5396_n6451.n177 AVSS 0.904589f
C6535 a_5396_n6451.t41 AVSS 0.323137f
C6536 a_5396_n6451.t18 AVSS 0.283144f
C6537 a_5396_n6451.t59 AVSS 0.24494f
C6538 a_5396_n6451.n178 AVSS 0.696106f
C6539 a_5396_n6451.t6 AVSS 0.242843f
C6540 a_5396_n6451.n179 AVSS 0.630724f
C6541 a_5396_n6451.t12 AVSS 0.283144f
C6542 a_5396_n6451.n180 AVSS 0.557056f
C6543 a_5396_n6451.t37 AVSS 0.242843f
C6544 a_5396_n6451.n181 AVSS 0.7005f
C6545 a_5396_n6451.t55 AVSS 0.244871f
C6546 a_5396_n6451.n182 AVSS 0.706241f
C6547 a_5396_n6451.t20 AVSS 0.283144f
C6548 a_5396_n6451.n183 AVSS 0.457093f
C6549 a_5396_n6451.n184 AVSS 0.160888f
C6550 a_5396_n6451.n185 AVSS 2.13459f
C6551 a_5396_n6451.n186 AVSS 2.37139f
C6552 a_5396_n6451.n187 AVSS 0.904589f
C6553 a_5396_n6451.t11 AVSS 0.323137f
C6554 a_5396_n6451.t39 AVSS 0.283144f
C6555 a_5396_n6451.t23 AVSS 0.24494f
C6556 a_5396_n6451.n188 AVSS 0.696106f
C6557 a_5396_n6451.t61 AVSS 0.242843f
C6558 a_5396_n6451.n189 AVSS 0.630724f
C6559 a_5396_n6451.n190 AVSS 0.815612f
C6560 a_5396_n6451.t56 AVSS 0.327688f
C6561 a_5396_n6451.t24 AVSS 0.283144f
C6562 a_5396_n6451.t66 AVSS 0.32522f
C6563 a_5396_n6451.t0 AVSS 0.278781f
C6564 a_5396_n6451.t64 AVSS 0.239195f
C6565 a_5396_n6451.n191 AVSS 0.715172f
C6566 a_5396_n6451.t65 AVSS 0.322023f
C6567 a_5396_n6451.n192 AVSS 1.2883f
C6568 a_5396_n6451.t1 AVSS 2.5812f
C6569 a_5396_n6451.t4 AVSS 0.550459f
C6570 a_5396_n6451.n193 AVSS 3.8859f
C6571 a_5396_n6451.t2 AVSS 0.783475f
C6572 a_5396_n6451.t63 AVSS 1.92091f
C6573 a_5396_n6451.t3 AVSS 0.322411f
C6574 a_5396_n6451.n194 AVSS 0.664255f
C6575 a_5396_n6451.n195 AVSS 2.8089f
C6576 a_5396_n6451.n196 AVSS 4.57358f
C6577 a_5396_n6451.t15 AVSS 0.326177f
C6578 a_5396_n6451.t35 AVSS 0.282702f
C6579 a_5396_n6451.t57 AVSS 0.244443f
C6580 a_5396_n6451.t36 AVSS 0.244125f
C6581 a_5396_n6451.n197 AVSS 3.69122f
C6582 a_5396_n6451.n198 AVSS 0.160881f
C6583 a_5396_n6451.t48 AVSS 0.282702f
C6584 a_5396_n6451.t40 AVSS 0.244443f
C6585 a_5396_n6451.t43 AVSS 0.244443f
C6586 a_5396_n6451.t13 AVSS 0.282702f
C6587 a_5396_n6451.t27 AVSS 0.244443f
C6588 a_5396_n6451.t50 AVSS 0.244125f
C6589 a_5396_n6451.t22 AVSS 0.282702f
C6590 a_5396_n6451.t32 AVSS 0.326614f
C6591 a_5396_n6451.n199 AVSS 0.160881f
C6592 a_5396_n6451.n200 AVSS 3.72221f
C6593 a_5396_n6451.t54 AVSS 1.08015f
C6594 a_5396_n6451.t47 AVSS 3.04535f
C6595 a_5396_n6451.t21 AVSS 1.86414f
C6596 a_5396_n6451.t9 AVSS 0.392888f
C6597 a_5396_n6451.t10 AVSS 1.21583f
C6598 a_5396_n6451.n201 AVSS 2.7314f
C6599 a_5396_n6451.n202 AVSS 2.11666f
C6600 a_5396_n6451.n203 AVSS 0.160888f
C6601 a_5396_n6451.t34 AVSS 0.242843f
C6602 a_5396_n6451.n204 AVSS 0.630724f
C6603 a_5396_n6451.t42 AVSS 0.24494f
C6604 a_5396_n6451.n205 AVSS 0.696106f
C6605 a_5396_n6451.t51 AVSS 0.283144f
C6606 a_5396_n6451.n206 AVSS 0.557056f
C6607 a_5396_n6451.t45 AVSS 0.242843f
C6608 a_5396_n6451.n207 AVSS 0.7005f
C6609 a_5396_n6451.t29 AVSS 0.244871f
C6610 a_5396_n6451.n208 AVSS 0.706241f
C6611 a_5396_n6451.t7 AVSS 0.283144f
C6612 a_5396_n6451.n209 AVSS 0.457093f
C6613 a_5396_n6451.n210 AVSS 0.160888f
C6614 a_5396_n6451.n211 AVSS 2.11666f
C6615 a_5396_n6451.t62 AVSS 0.326177f
C6616 a_5396_n6451.t53 AVSS 0.282702f
C6617 a_5396_n6451.t60 AVSS 0.244443f
C6618 a_5396_n6451.t58 AVSS 0.244125f
C6619 a_5396_n6451.t44 AVSS 0.282702f
C6620 a_5396_n6451.t33 AVSS 0.244443f
C6621 a_5396_n6451.t38 AVSS 0.244443f
C6622 a_5396_n6451.t26 AVSS 0.282702f
C6623 a_5396_n6451.t49 AVSS 0.244443f
C6624 a_5396_n6451.t46 AVSS 0.244125f
C6625 a_5396_n6451.t14 AVSS 0.282702f
C6626 a_5396_n6451.t19 AVSS 0.326614f
C6627 a_5396_n6451.n212 AVSS 0.160881f
C6628 a_5396_n6451.n213 AVSS 0.160881f
C6629 a_5396_n6451.n214 AVSS 2.35461f
C6630 a_5396_n6451.t25 AVSS 1.86414f
C6631 a_5396_n6451.t31 AVSS 0.392888f
C6632 a_5396_n6451.t30 AVSS 1.21583f
C6633 a_5396_n6451.n215 AVSS 2.7314f
C6634 a_5396_n6451.t28 AVSS 0.283144f
C6635 a_5396_n6451.n216 AVSS 0.815606f
C6636 a_5396_n6451.t5 AVSS 0.327695f
C6637 AVDD.t1187 AVSS 0.089409f
C6638 AVDD.t431 AVSS 0.089409f
C6639 AVDD.n0 AVSS 0.741323f
C6640 AVDD.t954 AVSS 0.045717f
C6641 AVDD.t416 AVSS 0.045717f
C6642 AVDD.t415 AVSS 0.089409f
C6643 AVDD.t320 AVSS 0.089409f
C6644 AVDD.t855 AVSS 0.045717f
C6645 AVDD.t321 AVSS 0.045717f
C6646 AVDD.n1 AVSS 0.378581f
C6647 AVDD.t924 AVSS 0.045717f
C6648 AVDD.t392 AVSS 0.045717f
C6649 AVDD.n2 AVSS 0.956364f
C6650 AVDD.n3 AVSS 0.374271f
C6651 AVDD.n4 AVSS 0.378609f
C6652 AVDD.n5 AVSS 16.0886f
C6653 AVDD.n6 AVSS 0.375467f
C6654 AVDD.n7 AVSS 0.375467f
C6655 AVDD.t70 AVSS 12.2951f
C6656 AVDD.n8 AVSS 0.374271f
C6657 AVDD.n9 AVSS 0.378609f
C6658 AVDD.t1060 AVSS 0.045717f
C6659 AVDD.t1070 AVSS 0.045717f
C6660 AVDD.n10 AVSS 0.872745f
C6661 AVDD.n11 AVSS 0.378581f
C6662 AVDD.t1066 AVSS 0.045717f
C6663 AVDD.t1090 AVSS 0.045717f
C6664 AVDD.t1089 AVSS 0.089409f
C6665 AVDD.t261 AVSS 0.089409f
C6666 AVDD.t760 AVSS 0.045717f
C6667 AVDD.t262 AVSS 0.045717f
C6668 AVDD.t314 AVSS 0.089409f
C6669 AVDD.t849 AVSS 0.045717f
C6670 AVDD.t315 AVSS 0.045717f
C6671 AVDD.n12 AVSS 0.301403f
C6672 AVDD.n13 AVSS 0.301403f
C6673 AVDD.t1226 AVSS 0.045717f
C6674 AVDD.t726 AVSS 0.045717f
C6675 AVDD.t725 AVSS 0.089409f
C6676 AVDD.t669 AVSS 0.045717f
C6677 AVDD.t129 AVSS 0.045717f
C6678 AVDD.t128 AVSS 0.089409f
C6679 AVDD.t266 AVSS 0.089409f
C6680 AVDD.t794 AVSS 0.045717f
C6681 AVDD.t267 AVSS 0.045717f
C6682 AVDD.n14 AVSS 0.378581f
C6683 AVDD.t782 AVSS 0.045717f
C6684 AVDD.t248 AVSS 0.045717f
C6685 AVDD.t247 AVSS 0.089409f
C6686 AVDD.t353 AVSS 0.089409f
C6687 AVDD.t890 AVSS 0.045717f
C6688 AVDD.t354 AVSS 0.045717f
C6689 AVDD.t1119 AVSS 0.089409f
C6690 AVDD.t371 AVSS 0.045717f
C6691 AVDD.t1120 AVSS 0.045717f
C6692 AVDD.n15 AVSS 0.153168f
C6693 AVDD.t1073 AVSS 0.089409f
C6694 AVDD.n16 AVSS 0.173626f
C6695 AVDD.t572 AVSS 0.021426f
C6696 AVDD.t170 AVSS 0.089409f
C6697 AVDD.n17 AVSS 0.173626f
C6698 AVDD.t184 AVSS 0.033572f
C6699 AVDD.t355 AVSS 0.089409f
C6700 AVDD.n18 AVSS 0.173626f
C6701 AVDD.t632 AVSS 0.021426f
C6702 AVDD.t631 AVSS 0.089409f
C6703 AVDD.n19 AVSS 0.110794f
C6704 AVDD.n20 AVSS 0.378581f
C6705 AVDD.t294 AVSS 13.1202f
C6706 AVDD.t141 AVSS 10.1876f
C6707 AVDD.t136 AVSS 10.1876f
C6708 AVDD.t153 AVSS 12.609f
C6709 AVDD.t5 AVSS 12.322001f
C6710 AVDD.n21 AVSS 0.378609f
C6711 AVDD.t98 AVSS 5.3808f
C6712 AVDD.n22 AVSS 0.374271f
C6713 AVDD.n23 AVSS 0.378581f
C6714 AVDD.n24 AVSS 0.26267f
C6715 AVDD.t1227 AVSS 0.089409f
C6716 AVDD.n25 AVSS 0.021426f
C6717 AVDD.t375 AVSS 0.089409f
C6718 AVDD.t1023 AVSS 0.089409f
C6719 AVDD.n26 AVSS 0.342362f
C6720 AVDD.t610 AVSS 0.021426f
C6721 AVDD.t376 AVSS 0.033572f
C6722 AVDD.t341 AVSS 0.033572f
C6723 AVDD.t340 AVSS 0.089409f
C6724 AVDD.t987 AVSS 0.089409f
C6725 AVDD.n27 AVSS 0.342362f
C6726 AVDD.t1242 AVSS 0.021426f
C6727 AVDD.n28 AVSS 0.021426f
C6728 AVDD.t617 AVSS 0.089409f
C6729 AVDD.t618 AVSS 0.021426f
C6730 AVDD.n29 AVSS 0.021426f
C6731 AVDD.t188 AVSS 0.089409f
C6732 AVDD.t852 AVSS 0.089409f
C6733 AVDD.n30 AVSS 0.342362f
C6734 AVDD.t1112 AVSS 0.033572f
C6735 AVDD.t189 AVSS 0.021426f
C6736 AVDD.n31 AVSS 0.021426f
C6737 AVDD.t465 AVSS 0.089409f
C6738 AVDD.t466 AVSS 0.033572f
C6739 AVDD.n32 AVSS 0.301403f
C6740 AVDD.t1236 AVSS 0.045717f
C6741 AVDD.t49 AVSS 0.045717f
C6742 AVDD.n33 AVSS 0.446747f
C6743 AVDD.t606 AVSS 0.045717f
C6744 AVDD.t720 AVSS 0.045717f
C6745 AVDD.t719 AVSS 0.089409f
C6746 AVDD.t1100 AVSS 0.045717f
C6747 AVDD.t1206 AVSS 0.045717f
C6748 AVDD.t1205 AVSS 0.089409f
C6749 AVDD.t1095 AVSS 0.089409f
C6750 AVDD.t1000 AVSS 0.045717f
C6751 AVDD.t1096 AVSS 0.045717f
C6752 AVDD.t882 AVSS 0.045717f
C6753 AVDD.t458 AVSS 0.045717f
C6754 AVDD.n34 AVSS 0.587661f
C6755 AVDD.n35 AVSS 0.374271f
C6756 AVDD.n36 AVSS 0.378609f
C6757 AVDD.t252 AVSS 12.609f
C6758 AVDD.t0 AVSS 12.609f
C6759 AVDD.t53 AVSS 10.1876f
C6760 AVDD.t30 AVSS 10.1876f
C6761 AVDD.t335 AVSS 13.1202f
C6762 AVDD.t16 AVSS 12.2951f
C6763 AVDD.n37 AVSS 5.56016f
C6764 AVDD.n38 AVSS 0.375467f
C6765 AVDD.t8 AVSS 8.42992f
C6766 AVDD.n39 AVSS 0.375467f
C6767 AVDD.n40 AVSS 0.374271f
C6768 AVDD.n41 AVSS 0.378609f
C6769 AVDD.n42 AVSS 0.148966f
C6770 AVDD.n43 AVSS 0.068966f
C6771 AVDD.t948 AVSS 0.021426f
C6772 AVDD.t947 AVSS 0.089409f
C6773 AVDD.n44 AVSS 0.169461f
C6774 AVDD.t1207 AVSS 0.089409f
C6775 AVDD.n45 AVSS 0.077127f
C6776 AVDD.n46 AVSS 0.379771f
C6777 AVDD.t1386 AVSS 0.010713f
C6778 AVDD.t1678 AVSS 0.010713f
C6779 AVDD.n47 AVSS 0.058856f
C6780 AVDD.t1297 AVSS 0.010713f
C6781 AVDD.t1294 AVSS 0.010713f
C6782 AVDD.n48 AVSS 0.039303f
C6783 AVDD.n49 AVSS 0.193299f
C6784 AVDD.t1402 AVSS 0.010713f
C6785 AVDD.t1446 AVSS 0.010713f
C6786 AVDD.n50 AVSS 0.039303f
C6787 AVDD.n51 AVSS 0.137092f
C6788 AVDD.t1433 AVSS 0.010713f
C6789 AVDD.t1491 AVSS 0.010713f
C6790 AVDD.n52 AVSS 0.039303f
C6791 AVDD.n53 AVSS 0.055061f
C6792 AVDD.n54 AVSS 0.055933f
C6793 AVDD.t818 AVSS 0.089409f
C6794 AVDD.n55 AVSS 0.077127f
C6795 AVDD.t63 AVSS 0.045717f
C6796 AVDD.n56 AVSS 0.37055f
C6797 AVDD.t869 AVSS 0.021426f
C6798 AVDD.t1247 AVSS 0.089409f
C6799 AVDD.n57 AVSS 0.169461f
C6800 AVDD.t996 AVSS 0.033572f
C6801 AVDD.t731 AVSS 0.089409f
C6802 AVDD.n58 AVSS 0.169461f
C6803 AVDD.t305 AVSS 0.021426f
C6804 AVDD.t342 AVSS 0.089409f
C6805 AVDD.n59 AVSS 0.169461f
C6806 AVDD.t585 AVSS 0.089409f
C6807 AVDD.n60 AVSS 0.169461f
C6808 AVDD.t146 AVSS 0.021426f
C6809 AVDD.t737 AVSS 0.089409f
C6810 AVDD.n61 AVSS 0.169461f
C6811 AVDD.t311 AVSS 0.033572f
C6812 AVDD.t310 AVSS 0.089409f
C6813 AVDD.n62 AVSS 0.149288f
C6814 AVDD.n63 AVSS 0.41016f
C6815 AVDD.t1167 AVSS 0.089409f
C6816 AVDD.n64 AVSS 0.149288f
C6817 AVDD.t642 AVSS 0.089409f
C6818 AVDD.n65 AVSS 0.169461f
C6819 AVDD.n66 AVSS 0.068966f
C6820 AVDD.t1008 AVSS 0.021426f
C6821 AVDD.t1007 AVSS 0.089409f
C6822 AVDD.n67 AVSS 0.169461f
C6823 AVDD.t138 AVSS 0.089409f
C6824 AVDD.n68 AVSS 0.077127f
C6825 AVDD.n69 AVSS 0.429161f
C6826 AVDD.t1527 AVSS 0.010713f
C6827 AVDD.t1339 AVSS 0.010713f
C6828 AVDD.n70 AVSS 0.058856f
C6829 AVDD.t1309 AVSS 0.010713f
C6830 AVDD.t1614 AVSS 0.010713f
C6831 AVDD.n71 AVSS 0.039303f
C6832 AVDD.n72 AVSS 0.193299f
C6833 AVDD.t1370 AVSS 0.010713f
C6834 AVDD.t1625 AVSS 0.010713f
C6835 AVDD.n73 AVSS 0.039303f
C6836 AVDD.n74 AVSS 0.137092f
C6837 AVDD.t1531 AVSS 0.010713f
C6838 AVDD.t1365 AVSS 0.010713f
C6839 AVDD.n75 AVSS 0.039303f
C6840 AVDD.n76 AVSS 0.055061f
C6841 AVDD.n77 AVSS 0.055933f
C6842 AVDD.t344 AVSS 0.089409f
C6843 AVDD.n78 AVSS 0.077127f
C6844 AVDD.n79 AVSS 0.585364f
C6845 AVDD.t780 AVSS 0.021426f
C6846 AVDD.t1161 AVSS 0.089409f
C6847 AVDD.n80 AVSS 0.169461f
C6848 AVDD.t307 AVSS 0.033572f
C6849 AVDD.t575 AVSS 0.089409f
C6850 AVDD.n81 AVSS 0.169461f
C6851 AVDD.t871 AVSS 0.021426f
C6852 AVDD.n82 AVSS 0.129712f
C6853 AVDD.n83 AVSS 0.375467f
C6854 AVDD.n84 AVSS 0.378581f
C6855 AVDD.t381 AVSS 12.322001f
C6856 AVDD.n85 AVSS 0.378609f
C6857 AVDD.n86 AVSS 0.378609f
C6858 AVDD.n87 AVSS 0.378609f
C6859 AVDD.n88 AVSS 0.378609f
C6860 AVDD.t88 AVSS 5.3808f
C6861 AVDD.n89 AVSS 0.374271f
C6862 AVDD.n90 AVSS 0.374271f
C6863 AVDD.n91 AVSS 0.375467f
C6864 AVDD.n92 AVSS 0.378581f
C6865 AVDD.n93 AVSS 0.26267f
C6866 AVDD.t87 AVSS 0.089409f
C6867 AVDD.n94 AVSS 0.021426f
C6868 AVDD.t1091 AVSS 0.089409f
C6869 AVDD.t455 AVSS 0.089409f
C6870 AVDD.n95 AVSS 0.342362f
C6871 AVDD.t764 AVSS 0.021426f
C6872 AVDD.t1092 AVSS 0.033572f
C6873 AVDD.t847 AVSS 0.033572f
C6874 AVDD.t846 AVSS 0.089409f
C6875 AVDD.t192 AVSS 0.089409f
C6876 AVDD.n96 AVSS 0.342362f
C6877 AVDD.t1034 AVSS 0.021426f
C6878 AVDD.n97 AVSS 0.021426f
C6879 AVDD.t403 AVSS 0.089409f
C6880 AVDD.t404 AVSS 0.021426f
C6881 AVDD.n98 AVSS 0.021426f
C6882 AVDD.t1267 AVSS 0.089409f
C6883 AVDD.t660 AVSS 0.089409f
C6884 AVDD.n99 AVSS 0.342362f
C6885 AVDD.t242 AVSS 0.033572f
C6886 AVDD.t1268 AVSS 0.021426f
C6887 AVDD.n100 AVSS 0.021426f
C6888 AVDD.t885 AVSS 0.089409f
C6889 AVDD.t886 AVSS 0.033572f
C6890 AVDD.n101 AVSS 0.301403f
C6891 AVDD.t96 AVSS 0.045717f
C6892 AVDD.t958 AVSS 0.045717f
C6893 AVDD.n102 AVSS 0.446747f
C6894 AVDD.t754 AVSS 0.045717f
C6895 AVDD.t319 AVSS 0.045717f
C6896 AVDD.t318 AVSS 0.089409f
C6897 AVDD.t1238 AVSS 0.045717f
C6898 AVDD.t837 AVSS 0.045717f
C6899 AVDD.t836 AVSS 0.089409f
C6900 AVDD.t721 AVSS 0.089409f
C6901 AVDD.t1144 AVSS 0.045717f
C6902 AVDD.t722 AVSS 0.045717f
C6903 AVDD.t499 AVSS 0.045717f
C6904 AVDD.t1220 AVSS 0.045717f
C6905 AVDD.n103 AVSS 0.587661f
C6906 AVDD.n104 AVSS 0.374271f
C6907 AVDD.n105 AVSS 0.378609f
C6908 AVDD.t59 AVSS 12.609f
C6909 AVDD.t193 AVSS 12.609f
C6910 AVDD.t279 AVSS 10.1876f
C6911 AVDD.t291 AVSS 10.1876f
C6912 AVDD.t241 AVSS 13.1202f
C6913 AVDD.t79 AVSS 12.2951f
C6914 AVDD.n106 AVSS 5.56016f
C6915 AVDD.n107 AVSS 0.375467f
C6916 AVDD.t56 AVSS 12.2951f
C6917 AVDD.n108 AVSS 0.375467f
C6918 AVDD.n109 AVSS 0.374271f
C6919 AVDD.n110 AVSS 0.139176f
C6920 AVDD.t178 AVSS 13.1202f
C6921 AVDD.t148 AVSS 10.1876f
C6922 AVDD.t111 AVSS 10.1876f
C6923 AVDD.t226 AVSS 12.609f
C6924 AVDD.t200 AVSS 12.322001f
C6925 AVDD.n111 AVSS 0.378609f
C6926 AVDD.n112 AVSS 0.378609f
C6927 AVDD.t114 AVSS 12.2951f
C6928 AVDD.t22 AVSS 13.1202f
C6929 AVDD.t119 AVSS 10.1876f
C6930 AVDD.t399 AVSS 10.1876f
C6931 AVDD.t338 AVSS 12.609f
C6932 AVDD.t156 AVSS 12.609f
C6933 AVDD.t175 AVSS 5.3808f
C6934 AVDD.n113 AVSS 0.374271f
C6935 AVDD.n114 AVSS 0.462621f
C6936 AVDD.t235 AVSS 0.089409f
C6937 AVDD.n115 AVSS 0.021426f
C6938 AVDD.t160 AVSS 0.089409f
C6939 AVDD.t155 AVSS 0.089409f
C6940 AVDD.n116 AVSS 0.55425f
C6941 AVDD.t473 AVSS 0.089409f
C6942 AVDD.t461 AVSS 0.089409f
C6943 AVDD.n117 AVSS 0.55425f
C6944 AVDD.t474 AVSS 0.033572f
C6945 AVDD.t535 AVSS 0.021426f
C6946 AVDD.t540 AVSS 0.089409f
C6947 AVDD.t534 AVSS 0.089409f
C6948 AVDD.n118 AVSS 0.55425f
C6949 AVDD.t173 AVSS 0.021426f
C6950 AVDD.t172 AVSS 0.089409f
C6951 AVDD.t164 AVSS 0.089409f
C6952 AVDD.n119 AVSS 0.55425f
C6953 AVDD.t244 AVSS 0.033572f
C6954 AVDD.t249 AVSS 0.089409f
C6955 AVDD.t243 AVSS 0.089409f
C6956 AVDD.n120 AVSS 0.55425f
C6957 AVDD.t975 AVSS 0.089409f
C6958 AVDD.t967 AVSS 0.089409f
C6959 AVDD.n121 AVSS 0.55425f
C6960 AVDD.t976 AVSS 0.045717f
C6961 AVDD.t1219 AVSS 0.089409f
C6962 AVDD.t498 AVSS 0.089409f
C6963 AVDD.n122 AVSS 0.445699f
C6964 AVDD.t1115 AVSS 0.089409f
C6965 AVDD.t389 AVSS 0.089409f
C6966 AVDD.n123 AVSS 0.445699f
C6967 AVDD.t390 AVSS 0.045717f
C6968 AVDD.t1116 AVSS 0.045717f
C6969 AVDD.n124 AVSS 0.743554f
C6970 AVDD.t198 AVSS 0.045717f
C6971 AVDD.t930 AVSS 0.045717f
C6972 AVDD.n125 AVSS 0.743554f
C6973 AVDD.t409 AVSS 0.089409f
C6974 AVDD.t407 AVSS 0.089409f
C6975 AVDD.n126 AVSS 0.55425f
C6976 AVDD.t410 AVSS 0.045717f
C6977 AVDD.t1155 AVSS 0.089409f
C6978 AVDD.t1147 AVSS 0.089409f
C6979 AVDD.n127 AVSS 0.55425f
C6980 AVDD.t1156 AVSS 0.033572f
C6981 AVDD.t786 AVSS 0.021426f
C6982 AVDD.t787 AVSS 0.089409f
C6983 AVDD.t785 AVSS 0.089409f
C6984 AVDD.n128 AVSS 0.55425f
C6985 AVDD.t865 AVSS 0.021426f
C6986 AVDD.t864 AVSS 0.089409f
C6987 AVDD.t856 AVSS 0.089409f
C6988 AVDD.n129 AVSS 0.55425f
C6989 AVDD.t460 AVSS 0.033572f
C6990 AVDD.t467 AVSS 0.089409f
C6991 AVDD.t459 AVSS 0.089409f
C6992 AVDD.n130 AVSS 0.55425f
C6993 AVDD.t860 AVSS 0.089409f
C6994 AVDD.t858 AVSS 0.089409f
C6995 AVDD.n131 AVSS 0.55425f
C6996 AVDD.t861 AVSS 0.033572f
C6997 AVDD.t908 AVSS 0.021426f
C6998 AVDD.t913 AVSS 0.089409f
C6999 AVDD.t907 AVSS 0.089409f
C7000 AVDD.n132 AVSS 0.33675f
C7001 AVDD.t539 AVSS 0.033572f
C7002 AVDD.t538 AVSS 0.089409f
C7003 AVDD.t530 AVSS 0.089409f
C7004 AVDD.n133 AVSS 0.55425f
C7005 AVDD.n134 AVSS 0.24512f
C7006 AVDD.t1229 AVSS 0.089409f
C7007 AVDD.t1223 AVSS 0.089409f
C7008 AVDD.n135 AVSS 0.55425f
C7009 AVDD.t1230 AVSS 0.033572f
C7010 AVDD.t1270 AVSS 0.021426f
C7011 AVDD.t1273 AVSS 0.089409f
C7012 AVDD.t1269 AVSS 0.089409f
C7013 AVDD.n136 AVSS 0.55425f
C7014 AVDD.t772 AVSS 0.021426f
C7015 AVDD.t771 AVSS 0.089409f
C7016 AVDD.t767 AVSS 0.089409f
C7017 AVDD.n137 AVSS 0.55425f
C7018 AVDD.t821 AVSS 0.033572f
C7019 AVDD.t828 AVSS 0.089409f
C7020 AVDD.t820 AVSS 0.089409f
C7021 AVDD.n138 AVSS 0.55425f
C7022 AVDD.t597 AVSS 0.089409f
C7023 AVDD.t591 AVSS 0.089409f
C7024 AVDD.n139 AVSS 0.411839f
C7025 AVDD.t598 AVSS 0.045717f
C7026 AVDD.n140 AVSS 0.241042f
C7027 AVDD.n141 AVSS 0.137622f
C7028 AVDD.t826 AVSS 0.089409f
C7029 AVDD.n142 AVSS 0.149288f
C7030 AVDD.t537 AVSS 0.021426f
C7031 AVDD.n143 AVSS 0.413506f
C7032 AVDD.t1358 AVSS 0.082269f
C7033 AVDD.t1633 AVSS 0.010713f
C7034 AVDD.t1545 AVSS 0.010713f
C7035 AVDD.n144 AVSS 0.042824f
C7036 AVDD.n145 AVSS 0.289878f
C7037 AVDD.t933 AVSS 0.089409f
C7038 AVDD.n146 AVSS 0.149288f
C7039 AVDD.t652 AVSS 0.089409f
C7040 AVDD.n147 AVSS 0.169461f
C7041 AVDD.n148 AVSS 0.148966f
C7042 AVDD.t934 AVSS 0.033572f
C7043 AVDD.t112 AVSS 0.021426f
C7044 AVDD.t1107 AVSS 0.089409f
C7045 AVDD.n149 AVSS 0.169461f
C7046 AVDD.t1075 AVSS 0.089409f
C7047 AVDD.n150 AVSS 0.169461f
C7048 AVDD.t671 AVSS 0.021426f
C7049 AVDD.t383 AVSS 0.089409f
C7050 AVDD.n151 AVSS 0.169461f
C7051 AVDD.t421 AVSS 0.089409f
C7052 AVDD.n152 AVSS 0.169461f
C7053 AVDD.t1264 AVSS 0.021426f
C7054 AVDD.n153 AVSS 0.021426f
C7055 AVDD.n154 AVSS 0.137456f
C7056 AVDD.t1263 AVSS 0.089409f
C7057 AVDD.n155 AVSS 0.169461f
C7058 AVDD.n156 AVSS 0.137456f
C7059 AVDD.n157 AVSS 0.021426f
C7060 AVDD.t422 AVSS 0.033572f
C7061 AVDD.n158 AVSS 0.144368f
C7062 AVDD.n159 AVSS 0.144368f
C7063 AVDD.t384 AVSS 0.033572f
C7064 AVDD.n160 AVSS 0.021426f
C7065 AVDD.n161 AVSS 0.137456f
C7066 AVDD.t670 AVSS 0.089409f
C7067 AVDD.n162 AVSS 0.108477f
C7068 AVDD.n163 AVSS 0.068728f
C7069 AVDD.n164 AVSS 0.129712f
C7070 AVDD.n165 AVSS 0.021426f
C7071 AVDD.t1076 AVSS 0.033572f
C7072 AVDD.n166 AVSS 0.144368f
C7073 AVDD.n167 AVSS 0.144368f
C7074 AVDD.t1108 AVSS 0.033572f
C7075 AVDD.n168 AVSS 0.021426f
C7076 AVDD.n169 AVSS 0.137456f
C7077 AVDD.t110 AVSS 0.089409f
C7078 AVDD.n170 AVSS 0.169461f
C7079 AVDD.n171 AVSS 0.137456f
C7080 AVDD.n172 AVSS 0.021426f
C7081 AVDD.t653 AVSS 0.021426f
C7082 AVDD.n173 AVSS 0.021426f
C7083 AVDD.n174 AVSS 0.117034f
C7084 AVDD.n175 AVSS 0.06773f
C7085 AVDD.n176 AVSS 0.453573f
C7086 AVDD.n177 AVSS 0.006326f
C7087 AVDD.n178 AVSS 0.006326f
C7088 AVDD.n179 AVSS 0.128885f
C7089 AVDD.t1321 AVSS 0.010713f
C7090 AVDD.t1554 AVSS 0.010713f
C7091 AVDD.n180 AVSS 0.03213f
C7092 AVDD.t1328 AVSS 0.010713f
C7093 AVDD.t1530 AVSS 0.010713f
C7094 AVDD.n181 AVSS 0.024902f
C7095 AVDD.n182 AVSS 0.103112f
C7096 AVDD.t1519 AVSS 0.010713f
C7097 AVDD.t1351 AVSS 0.010713f
C7098 AVDD.n183 AVSS 0.03213f
C7099 AVDD.t1496 AVSS 0.010713f
C7100 AVDD.t1322 AVSS 0.010713f
C7101 AVDD.n184 AVSS 0.024902f
C7102 AVDD.n185 AVSS 0.073953f
C7103 AVDD.n186 AVSS 0.148993f
C7104 AVDD.t1340 AVSS 0.010713f
C7105 AVDD.t1307 AVSS 0.010713f
C7106 AVDD.n187 AVSS 0.03213f
C7107 AVDD.t1521 AVSS 0.010713f
C7108 AVDD.t1378 AVSS 0.010713f
C7109 AVDD.n188 AVSS 0.024902f
C7110 AVDD.n189 AVSS 0.073953f
C7111 AVDD.n190 AVSS 0.115393f
C7112 AVDD.t1330 AVSS 0.010713f
C7113 AVDD.t1637 AVSS 0.010713f
C7114 AVDD.n191 AVSS 0.03213f
C7115 AVDD.t1558 AVSS 0.010713f
C7116 AVDD.t1344 AVSS 0.010713f
C7117 AVDD.n192 AVSS 0.024902f
C7118 AVDD.n193 AVSS 0.073953f
C7119 AVDD.n194 AVSS 0.030661f
C7120 AVDD.n195 AVSS 0.006326f
C7121 AVDD.n196 AVSS 0.006326f
C7122 AVDD.t1537 AVSS 0.027903f
C7123 AVDD.n197 AVSS 0.038333f
C7124 AVDD.n198 AVSS 0.014056f
C7125 AVDD.n199 AVSS 0.025752f
C7126 AVDD.n200 AVSS 0.025734f
C7127 AVDD.t1630 AVSS 0.010713f
C7128 AVDD.t1497 AVSS 0.010713f
C7129 AVDD.n201 AVSS 0.026809f
C7130 AVDD.n202 AVSS 0.027694f
C7131 AVDD.n203 AVSS 0.014056f
C7132 AVDD.n204 AVSS 0.149628f
C7133 AVDD.n205 AVSS 0.006326f
C7134 AVDD.t1333 AVSS 0.027903f
C7135 AVDD.n206 AVSS 0.038333f
C7136 AVDD.t1352 AVSS 0.010713f
C7137 AVDD.t1361 AVSS 0.010713f
C7138 AVDD.n207 AVSS 0.092646f
C7139 AVDD.n208 AVSS 0.199269f
C7140 AVDD.n209 AVSS 0.014056f
C7141 AVDD.n210 AVSS 0.054035f
C7142 AVDD.n211 AVSS 0.283675f
C7143 AVDD.n212 AVSS 0.632147f
C7144 AVDD.n213 AVSS 0.0901f
C7145 AVDD.t1619 AVSS 0.010713f
C7146 AVDD.t1533 AVSS 0.010713f
C7147 AVDD.n214 AVSS 0.03213f
C7148 AVDD.t1636 AVSS 0.010713f
C7149 AVDD.t1316 AVSS 0.010713f
C7150 AVDD.n215 AVSS 0.024902f
C7151 AVDD.n216 AVSS 0.073953f
C7152 AVDD.n217 AVSS 0.113804f
C7153 AVDD.t1539 AVSS 0.010713f
C7154 AVDD.t1371 AVSS 0.010713f
C7155 AVDD.n218 AVSS 0.03213f
C7156 AVDD.t1529 AVSS 0.010713f
C7157 AVDD.t1624 AVSS 0.010713f
C7158 AVDD.n219 AVSS 0.024902f
C7159 AVDD.n220 AVSS 0.073953f
C7160 AVDD.n221 AVSS 0.115396f
C7161 AVDD.t1549 AVSS 0.010713f
C7162 AVDD.t1360 AVSS 0.010713f
C7163 AVDD.n222 AVSS 0.03213f
C7164 AVDD.t1366 AVSS 0.010713f
C7165 AVDD.t1304 AVSS 0.010713f
C7166 AVDD.n223 AVSS 0.024902f
C7167 AVDD.n224 AVSS 0.073953f
C7168 AVDD.n225 AVSS 0.115393f
C7169 AVDD.t1613 AVSS 0.010713f
C7170 AVDD.t1510 AVSS 0.010713f
C7171 AVDD.n226 AVSS 0.03213f
C7172 AVDD.t1626 AVSS 0.010713f
C7173 AVDD.t1639 AVSS 0.010713f
C7174 AVDD.n227 AVSS 0.024902f
C7175 AVDD.n228 AVSS 0.073953f
C7176 AVDD.n229 AVSS 0.06419f
C7177 AVDD.n230 AVSS 0.715915f
C7178 AVDD.t1515 AVSS 0.082269f
C7179 AVDD.t1364 AVSS 0.010713f
C7180 AVDD.t1616 AVSS 0.010713f
C7181 AVDD.n231 AVSS 0.042824f
C7182 AVDD.n232 AVSS 0.289878f
C7183 AVDD.n233 AVSS 0.203305f
C7184 AVDD.t1631 AVSS 0.04243f
C7185 AVDD.n234 AVSS 0.202316f
C7186 AVDD.t1341 AVSS 0.010713f
C7187 AVDD.t1327 AVSS 0.010713f
C7188 AVDD.n235 AVSS 0.042824f
C7189 AVDD.n236 AVSS 0.156341f
C7190 AVDD.n237 AVSS 0.519769f
C7191 AVDD.n238 AVSS 0.447556f
C7192 AVDD.n239 AVSS 0.081607f
C7193 AVDD.t1318 AVSS 0.027903f
C7194 AVDD.n240 AVSS 0.038333f
C7195 AVDD.n241 AVSS 0.014056f
C7196 AVDD.n242 AVSS 0.025752f
C7197 AVDD.n243 AVSS 0.025734f
C7198 AVDD.t1500 AVSS 0.010713f
C7199 AVDD.t1536 AVSS 0.010713f
C7200 AVDD.n244 AVSS 0.026809f
C7201 AVDD.n245 AVSS 0.027694f
C7202 AVDD.n246 AVSS 0.014056f
C7203 AVDD.n247 AVSS 0.149628f
C7204 AVDD.n248 AVSS 0.006326f
C7205 AVDD.t1611 AVSS 0.027903f
C7206 AVDD.n249 AVSS 0.038333f
C7207 AVDD.t1524 AVSS 0.010713f
C7208 AVDD.t1557 AVSS 0.010713f
C7209 AVDD.n250 AVSS 0.092646f
C7210 AVDD.n251 AVSS 0.199269f
C7211 AVDD.n252 AVSS 0.014056f
C7212 AVDD.n253 AVSS 0.054035f
C7213 AVDD.n254 AVSS 0.197145f
C7214 AVDD.n255 AVSS 0.406385f
C7215 AVDD.t1540 AVSS 0.010713f
C7216 AVDD.t1353 AVSS 0.010713f
C7217 AVDD.n256 AVSS 0.03213f
C7218 AVDD.t1528 AVSS 0.010713f
C7219 AVDD.t1342 AVSS 0.010713f
C7220 AVDD.n257 AVSS 0.024902f
C7221 AVDD.n258 AVSS 0.073953f
C7222 AVDD.n259 AVSS 0.06419f
C7223 AVDD.t1324 AVSS 0.010713f
C7224 AVDD.t1628 AVSS 0.010713f
C7225 AVDD.n260 AVSS 0.03213f
C7226 AVDD.t1312 AVSS 0.010713f
C7227 AVDD.t1617 AVSS 0.010713f
C7228 AVDD.n261 AVSS 0.024902f
C7229 AVDD.n262 AVSS 0.073953f
C7230 AVDD.n263 AVSS 0.115393f
C7231 AVDD.t1313 AVSS 0.010713f
C7232 AVDD.t1499 AVSS 0.010713f
C7233 AVDD.n264 AVSS 0.03213f
C7234 AVDD.t1306 AVSS 0.010713f
C7235 AVDD.t1627 AVSS 0.010713f
C7236 AVDD.n265 AVSS 0.024902f
C7237 AVDD.n266 AVSS 0.073953f
C7238 AVDD.n267 AVSS 0.115396f
C7239 AVDD.t1548 AVSS 0.010713f
C7240 AVDD.t1310 AVSS 0.010713f
C7241 AVDD.n268 AVSS 0.03213f
C7242 AVDD.t1538 AVSS 0.010713f
C7243 AVDD.t1369 AVSS 0.010713f
C7244 AVDD.n269 AVSS 0.024902f
C7245 AVDD.n270 AVSS 0.073953f
C7246 AVDD.n271 AVSS 0.113804f
C7247 AVDD.t1516 AVSS 0.010713f
C7248 AVDD.t1334 AVSS 0.010713f
C7249 AVDD.n272 AVSS 0.03213f
C7250 AVDD.t1507 AVSS 0.010713f
C7251 AVDD.t1323 AVSS 0.010713f
C7252 AVDD.n273 AVSS 0.024902f
C7253 AVDD.n274 AVSS 0.103112f
C7254 AVDD.t1367 AVSS 0.010713f
C7255 AVDD.t1620 AVSS 0.010713f
C7256 AVDD.n275 AVSS 0.03213f
C7257 AVDD.t1356 AVSS 0.010713f
C7258 AVDD.t1609 AVSS 0.010713f
C7259 AVDD.n276 AVSS 0.024902f
C7260 AVDD.n277 AVSS 0.073953f
C7261 AVDD.n278 AVSS 0.148993f
C7262 AVDD.t1605 AVSS 0.010713f
C7263 AVDD.t1503 AVSS 0.010713f
C7264 AVDD.n279 AVSS 0.03213f
C7265 AVDD.t1329 AVSS 0.010713f
C7266 AVDD.t1635 AVSS 0.010713f
C7267 AVDD.n280 AVSS 0.024902f
C7268 AVDD.n281 AVSS 0.073953f
C7269 AVDD.n282 AVSS 0.115393f
C7270 AVDD.t1525 AVSS 0.010713f
C7271 AVDD.t1561 AVSS 0.010713f
C7272 AVDD.n283 AVSS 0.03213f
C7273 AVDD.t1517 AVSS 0.010713f
C7274 AVDD.t1552 AVSS 0.010713f
C7275 AVDD.n284 AVSS 0.024902f
C7276 AVDD.n285 AVSS 0.073953f
C7277 AVDD.n286 AVSS 0.030661f
C7278 AVDD.n287 AVSS 0.0901f
C7279 AVDD.n288 AVSS 0.41016f
C7280 AVDD.n289 AVSS 0.368072f
C7281 AVDD.n290 AVSS 0.203305f
C7282 AVDD.t1555 AVSS 0.04243f
C7283 AVDD.n291 AVSS 0.202316f
C7284 AVDD.t1607 AVSS 0.010713f
C7285 AVDD.t1520 AVSS 0.010713f
C7286 AVDD.n292 AVSS 0.042824f
C7287 AVDD.n293 AVSS 0.156341f
C7288 AVDD.n294 AVSS 0.434267f
C7289 AVDD.n295 AVSS 0.06773f
C7290 AVDD.t223 AVSS 0.089409f
C7291 AVDD.n296 AVSS 0.169461f
C7292 AVDD.t1214 AVSS 0.033572f
C7293 AVDD.t1253 AVSS 0.089409f
C7294 AVDD.n297 AVSS 0.169461f
C7295 AVDD.n298 AVSS 0.021426f
C7296 AVDD.t1254 AVSS 0.033572f
C7297 AVDD.n299 AVSS 0.144368f
C7298 AVDD.n300 AVSS 0.144368f
C7299 AVDD.t1213 AVSS 0.089409f
C7300 AVDD.n301 AVSS 0.169461f
C7301 AVDD.n302 AVSS 0.137456f
C7302 AVDD.n303 AVSS 0.021426f
C7303 AVDD.t224 AVSS 0.021426f
C7304 AVDD.n304 AVSS 0.021426f
C7305 AVDD.n305 AVSS 0.137456f
C7306 AVDD.t536 AVSS 0.089409f
C7307 AVDD.n306 AVSS 0.169461f
C7308 AVDD.n307 AVSS 0.117034f
C7309 AVDD.n308 AVSS 0.021426f
C7310 AVDD.t827 AVSS 0.033572f
C7311 AVDD.n309 AVSS 0.182536f
C7312 AVDD.t1038 AVSS 0.045717f
C7313 AVDD.n310 AVSS 0.37868f
C7314 AVDD.t1037 AVSS 0.089409f
C7315 AVDD.n311 AVSS 0.398711f
C7316 AVDD.t297 AVSS 0.045717f
C7317 AVDD.n312 AVSS 0.387307f
C7318 AVDD.t296 AVSS 0.089409f
C7319 AVDD.n313 AVSS 0.225482f
C7320 AVDD.t158 AVSS 0.089409f
C7321 AVDD.n314 AVSS 0.225482f
C7322 AVDD.t159 AVSS 0.045717f
C7323 AVDD.n315 AVSS 0.178363f
C7324 AVDD.n316 AVSS 0.170808f
C7325 AVDD.n317 AVSS 0.287122f
C7326 AVDD.t260 AVSS 0.045717f
C7327 AVDD.n318 AVSS 0.297599f
C7328 AVDD.t259 AVSS 0.089409f
C7329 AVDD.n319 AVSS 0.225482f
C7330 AVDD.t427 AVSS 0.089409f
C7331 AVDD.n320 AVSS 0.225482f
C7332 AVDD.t428 AVSS 0.045717f
C7333 AVDD.n321 AVSS 0.376621f
C7334 AVDD.n322 AVSS 0.236716f
C7335 AVDD.t308 AVSS 0.089409f
C7336 AVDD.t309 AVSS 0.045717f
C7337 AVDD.t45 AVSS 0.033572f
C7338 AVDD.t43 AVSS 0.089409f
C7339 AVDD.t727 AVSS 0.089409f
C7340 AVDD.n323 AVSS 0.342362f
C7341 AVDD.t424 AVSS 0.021426f
C7342 AVDD.n324 AVSS 0.021426f
C7343 AVDD.t1057 AVSS 0.089409f
C7344 AVDD.t1058 AVSS 0.021426f
C7345 AVDD.n325 AVSS 0.021426f
C7346 AVDD.t777 AVSS 0.089409f
C7347 AVDD.t121 AVSS 0.089409f
C7348 AVDD.n326 AVSS 0.342362f
C7349 AVDD.t1128 AVSS 0.033572f
C7350 AVDD.t778 AVSS 0.021426f
C7351 AVDD.n327 AVSS 0.021426f
C7352 AVDD.t482 AVSS 0.089409f
C7353 AVDD.t483 AVSS 0.033572f
C7354 AVDD.t89 AVSS 0.021426f
C7355 AVDD.n328 AVSS 0.021426f
C7356 AVDD.t525 AVSS 0.033572f
C7357 AVDD.t524 AVSS 0.089409f
C7358 AVDD.t1171 AVSS 0.089409f
C7359 AVDD.n329 AVSS 0.342362f
C7360 AVDD.n330 AVSS 0.021426f
C7361 AVDD.t1172 AVSS 0.033572f
C7362 AVDD.n331 AVSS 0.292092f
C7363 AVDD.n332 AVSS 0.292092f
C7364 AVDD.t1127 AVSS 0.089409f
C7365 AVDD.n333 AVSS 0.342362f
C7366 AVDD.n334 AVSS 0.278352f
C7367 AVDD.n335 AVSS 0.021426f
C7368 AVDD.t123 AVSS 0.021426f
C7369 AVDD.n336 AVSS 0.021426f
C7370 AVDD.n337 AVSS 0.278352f
C7371 AVDD.t423 AVSS 0.089409f
C7372 AVDD.n338 AVSS 0.342362f
C7373 AVDD.n339 AVSS 0.278352f
C7374 AVDD.n340 AVSS 0.021426f
C7375 AVDD.t728 AVSS 0.033572f
C7376 AVDD.n341 AVSS 0.320025f
C7377 AVDD.t952 AVSS 0.045717f
C7378 AVDD.n342 AVSS 0.320025f
C7379 AVDD.t951 AVSS 0.089409f
C7380 AVDD.n343 AVSS 0.261503f
C7381 AVDD.n344 AVSS 0.68361f
C7382 AVDD.t823 AVSS 0.045717f
C7383 AVDD.n345 AVSS 0.376621f
C7384 AVDD.t822 AVSS 0.089409f
C7385 AVDD.n346 AVSS 0.225482f
C7386 AVDD.t710 AVSS 0.089409f
C7387 AVDD.n347 AVSS 0.225482f
C7388 AVDD.t711 AVSS 0.045717f
C7389 AVDD.n348 AVSS 0.27229f
C7390 AVDD.n349 AVSS 0.180541f
C7391 AVDD.n350 AVSS 0.195047f
C7392 AVDD.t125 AVSS 0.045717f
C7393 AVDD.n351 AVSS 0.284944f
C7394 AVDD.t124 AVSS 0.089409f
C7395 AVDD.n352 AVSS 0.225482f
C7396 AVDD.t1271 AVSS 0.089409f
C7397 AVDD.n353 AVSS 0.225482f
C7398 AVDD.t1272 AVSS 0.045717f
C7399 AVDD.n354 AVSS 0.376621f
C7400 AVDD.t1094 AVSS 0.045717f
C7401 AVDD.t998 AVSS 0.045717f
C7402 AVDD.n355 AVSS 0.195241f
C7403 AVDD.t101 AVSS 0.045717f
C7404 AVDD.n356 AVSS 0.27229f
C7405 AVDD.n357 AVSS 0.137577f
C7406 AVDD.t68 AVSS 0.045717f
C7407 AVDD.t203 AVSS 0.045717f
C7408 AVDD.t980 AVSS 0.045717f
C7409 AVDD.t749 AVSS 0.089409f
C7410 AVDD.n358 AVSS 0.173626f
C7411 AVDD.t446 AVSS 0.021426f
C7412 AVDD.t133 AVSS 0.089409f
C7413 AVDD.n359 AVSS 0.173626f
C7414 AVDD.t1160 AVSS 0.033572f
C7415 AVDD.t1189 AVSS 0.089409f
C7416 AVDD.n360 AVSS 0.173626f
C7417 AVDD.t792 AVSS 0.021426f
C7418 AVDD.t490 AVSS 0.089409f
C7419 AVDD.n361 AVSS 0.173626f
C7420 AVDD.t217 AVSS 0.089409f
C7421 AVDD.n362 AVSS 0.173626f
C7422 AVDD.t1062 AVSS 0.021426f
C7423 AVDD.t688 AVSS 0.089409f
C7424 AVDD.n363 AVSS 0.173626f
C7425 AVDD.t275 AVSS 0.033572f
C7426 AVDD.t872 AVSS 0.089409f
C7427 AVDD.n364 AVSS 0.173626f
C7428 AVDD.t580 AVSS 0.021426f
C7429 AVDD.t1277 AVSS 0.089409f
C7430 AVDD.n365 AVSS 0.173626f
C7431 AVDD.t1028 AVSS 0.033572f
C7432 AVDD.t1011 AVSS 0.089409f
C7433 AVDD.n366 AVSS 0.173626f
C7434 AVDD.t590 AVSS 0.021426f
C7435 AVDD.t316 AVSS 0.089409f
C7436 AVDD.n367 AVSS 0.173626f
C7437 AVDD.t359 AVSS 0.089409f
C7438 AVDD.n368 AVSS 0.173626f
C7439 AVDD.t1202 AVSS 0.021426f
C7440 AVDD.t943 AVSS 0.089409f
C7441 AVDD.n369 AVSS 0.173626f
C7442 AVDD.t51 AVSS 0.033572f
C7443 AVDD.t50 AVSS 0.089409f
C7444 AVDD.n370 AVSS 0.173626f
C7445 AVDD.n371 AVSS 0.141621f
C7446 AVDD.n372 AVSS 0.021426f
C7447 AVDD.t944 AVSS 0.021426f
C7448 AVDD.n373 AVSS 0.021426f
C7449 AVDD.n374 AVSS 0.141621f
C7450 AVDD.t1201 AVSS 0.089409f
C7451 AVDD.n375 AVSS 0.173626f
C7452 AVDD.n376 AVSS 0.141621f
C7453 AVDD.n377 AVSS 0.021426f
C7454 AVDD.t360 AVSS 0.033572f
C7455 AVDD.n378 AVSS 0.148431f
C7456 AVDD.n379 AVSS 0.148431f
C7457 AVDD.t317 AVSS 0.033572f
C7458 AVDD.n380 AVSS 0.021426f
C7459 AVDD.n381 AVSS 0.141621f
C7460 AVDD.t589 AVSS 0.089409f
C7461 AVDD.n382 AVSS 0.110794f
C7462 AVDD.n383 AVSS 0.07081f
C7463 AVDD.n384 AVSS 0.133642f
C7464 AVDD.n385 AVSS 0.021426f
C7465 AVDD.t1012 AVSS 0.033572f
C7466 AVDD.n386 AVSS 0.148431f
C7467 AVDD.n387 AVSS 0.148431f
C7468 AVDD.t1027 AVSS 0.089409f
C7469 AVDD.n388 AVSS 0.173626f
C7470 AVDD.n389 AVSS 0.141621f
C7471 AVDD.n390 AVSS 0.021426f
C7472 AVDD.t1278 AVSS 0.021426f
C7473 AVDD.n391 AVSS 0.021426f
C7474 AVDD.n392 AVSS 0.141621f
C7475 AVDD.t579 AVSS 0.089409f
C7476 AVDD.n393 AVSS 0.173626f
C7477 AVDD.n394 AVSS 0.141621f
C7478 AVDD.n395 AVSS 0.021426f
C7479 AVDD.t873 AVSS 0.033572f
C7480 AVDD.n396 AVSS 0.153168f
C7481 AVDD.t434 AVSS 0.033572f
C7482 AVDD.t433 AVSS 0.089409f
C7483 AVDD.t1279 AVSS 0.089409f
C7484 AVDD.n397 AVSS 0.342362f
C7485 AVDD.t1030 AVSS 0.021426f
C7486 AVDD.n398 AVSS 0.021426f
C7487 AVDD.t147 AVSS 0.089409f
C7488 AVDD.t149 AVSS 0.021426f
C7489 AVDD.n399 AVSS 0.021426f
C7490 AVDD.t915 AVSS 0.089409f
C7491 AVDD.t504 AVSS 0.089409f
C7492 AVDD.n400 AVSS 0.342362f
C7493 AVDD.t227 AVSS 0.033572f
C7494 AVDD.t916 AVSS 0.021426f
C7495 AVDD.n401 AVSS 0.021426f
C7496 AVDD.t629 AVSS 0.089409f
C7497 AVDD.t630 AVSS 0.033572f
C7498 AVDD.t612 AVSS 0.033572f
C7499 AVDD.t611 AVSS 0.089409f
C7500 AVDD.t199 AVSS 0.089409f
C7501 AVDD.n402 AVSS 0.342362f
C7502 AVDD.t1052 AVSS 0.021426f
C7503 AVDD.n403 AVSS 0.021426f
C7504 AVDD.t174 AVSS 0.089409f
C7505 AVDD.t176 AVSS 0.021426f
C7506 AVDD.n404 AVSS 0.021426f
C7507 AVDD.t1175 AVSS 0.089409f
C7508 AVDD.t795 AVSS 0.089409f
C7509 AVDD.n405 AVSS 0.342362f
C7510 AVDD.t1176 AVSS 0.033572f
C7511 AVDD.t1218 AVSS 0.033572f
C7512 AVDD.t1217 AVSS 0.089409f
C7513 AVDD.t838 AVSS 0.089409f
C7514 AVDD.n406 AVSS 0.342362f
C7515 AVDD.t400 AVSS 0.021426f
C7516 AVDD.n407 AVSS 0.021426f
C7517 AVDD.t814 AVSS 0.089409f
C7518 AVDD.t815 AVSS 0.021426f
C7519 AVDD.n408 AVSS 0.021426f
C7520 AVDD.t522 AVSS 0.089409f
C7521 AVDD.t118 AVSS 0.089409f
C7522 AVDD.n409 AVSS 0.342362f
C7523 AVDD.t558 AVSS 0.033572f
C7524 AVDD.t523 AVSS 0.021426f
C7525 AVDD.t950 AVSS 0.033572f
C7526 AVDD.n410 AVSS 0.021426f
C7527 AVDD.t949 AVSS 0.089409f
C7528 AVDD.t557 AVSS 0.089409f
C7529 AVDD.n411 AVSS 0.342362f
C7530 AVDD.n412 AVSS 0.278352f
C7531 AVDD.n413 AVSS 0.021426f
C7532 AVDD.t120 AVSS 0.021426f
C7533 AVDD.n414 AVSS 0.021426f
C7534 AVDD.n415 AVSS 0.278352f
C7535 AVDD.t398 AVSS 0.089409f
C7536 AVDD.n416 AVSS 0.342362f
C7537 AVDD.n417 AVSS 0.278352f
C7538 AVDD.n418 AVSS 0.021426f
C7539 AVDD.t839 AVSS 0.033572f
C7540 AVDD.n419 AVSS 0.292092f
C7541 AVDD.n420 AVSS 0.292092f
C7542 AVDD.t796 AVSS 0.033572f
C7543 AVDD.n421 AVSS 0.021426f
C7544 AVDD.n422 AVSS 0.278352f
C7545 AVDD.t1051 AVSS 0.089409f
C7546 AVDD.n423 AVSS 0.218868f
C7547 AVDD.n424 AVSS 0.139176f
C7548 AVDD.n425 AVSS 0.26267f
C7549 AVDD.n426 AVSS 0.021426f
C7550 AVDD.t201 AVSS 0.033572f
C7551 AVDD.n427 AVSS 0.292092f
C7552 AVDD.n428 AVSS 0.292092f
C7553 AVDD.t225 AVSS 0.089409f
C7554 AVDD.n429 AVSS 0.342362f
C7555 AVDD.n430 AVSS 0.278352f
C7556 AVDD.n431 AVSS 0.021426f
C7557 AVDD.t505 AVSS 0.021426f
C7558 AVDD.n432 AVSS 0.021426f
C7559 AVDD.n433 AVSS 0.278352f
C7560 AVDD.t1029 AVSS 0.089409f
C7561 AVDD.n434 AVSS 0.342362f
C7562 AVDD.n435 AVSS 0.278352f
C7563 AVDD.n436 AVSS 0.021426f
C7564 AVDD.t1280 AVSS 0.033572f
C7565 AVDD.n437 AVSS 0.301403f
C7566 AVDD.t929 AVSS 0.089409f
C7567 AVDD.t197 AVSS 0.089409f
C7568 AVDD.n438 AVSS 0.445699f
C7569 AVDD.t824 AVSS 0.089409f
C7570 AVDD.t55 AVSS 0.089409f
C7571 AVDD.n439 AVSS 0.445699f
C7572 AVDD.t57 AVSS 0.045717f
C7573 AVDD.t825 AVSS 0.045717f
C7574 AVDD.n440 AVSS 0.537731f
C7575 AVDD.n441 AVSS 0.378581f
C7576 AVDD.n442 AVSS 0.712338f
C7577 AVDD.t75 AVSS 0.045717f
C7578 AVDD.t843 AVSS 0.045717f
C7579 AVDD.n443 AVSS 0.587661f
C7580 AVDD.t842 AVSS 0.089409f
C7581 AVDD.t74 AVSS 0.089409f
C7582 AVDD.n444 AVSS 0.445699f
C7583 AVDD.t830 AVSS 0.089409f
C7584 AVDD.t546 AVSS 0.089409f
C7585 AVDD.n445 AVSS 0.445699f
C7586 AVDD.t547 AVSS 0.045717f
C7587 AVDD.t831 AVSS 0.045717f
C7588 AVDD.n446 AVSS 0.764636f
C7589 AVDD.t162 AVSS 0.089409f
C7590 AVDD.t603 AVSS 0.089409f
C7591 AVDD.n447 AVSS 0.787444f
C7592 AVDD.t604 AVSS 0.045717f
C7593 AVDD.t163 AVSS 0.045717f
C7594 AVDD.n448 AVSS 0.446747f
C7595 AVDD.t1139 AVSS 0.089409f
C7596 AVDD.t735 AVSS 0.089409f
C7597 AVDD.n449 AVSS 0.342362f
C7598 AVDD.t1140 AVSS 0.033572f
C7599 AVDD.t1164 AVSS 0.021426f
C7600 AVDD.t290 AVSS 0.089409f
C7601 AVDD.t1163 AVSS 0.089409f
C7602 AVDD.n450 AVSS 0.342362f
C7603 AVDD.t675 AVSS 0.021426f
C7604 AVDD.t674 AVSS 0.089409f
C7605 AVDD.t278 AVSS 0.089409f
C7606 AVDD.n451 AVSS 0.342362f
C7607 AVDD.t699 AVSS 0.033572f
C7608 AVDD.t1077 AVSS 0.089409f
C7609 AVDD.t698 AVSS 0.089409f
C7610 AVDD.n452 AVSS 0.342362f
C7611 AVDD.t58 AVSS 0.089409f
C7612 AVDD.t969 AVSS 0.089409f
C7613 AVDD.n453 AVSS 0.342362f
C7614 AVDD.t60 AVSS 0.033572f
C7615 AVDD.t1234 AVSS 0.021426f
C7616 AVDD.t363 AVSS 0.089409f
C7617 AVDD.t1233 AVSS 0.089409f
C7618 AVDD.n454 AVSS 0.218868f
C7619 AVDD.t804 AVSS 0.033572f
C7620 AVDD.t803 AVSS 0.089409f
C7621 AVDD.t380 AVSS 0.089409f
C7622 AVDD.n455 AVSS 0.342362f
C7623 AVDD.n456 AVSS 0.139176f
C7624 AVDD.t757 AVSS 0.089409f
C7625 AVDD.t346 AVSS 0.089409f
C7626 AVDD.n457 AVSS 0.342362f
C7627 AVDD.t758 AVSS 0.033572f
C7628 AVDD.t624 AVSS 0.021426f
C7629 AVDD.t1021 AVSS 0.089409f
C7630 AVDD.t623 AVSS 0.089409f
C7631 AVDD.n458 AVSS 0.342362f
C7632 AVDD.t20 AVSS 0.021426f
C7633 AVDD.t18 AVSS 0.089409f
C7634 AVDD.t939 AVSS 0.089409f
C7635 AVDD.n459 AVSS 0.342362f
C7636 AVDD.t1200 AVSS 0.033572f
C7637 AVDD.t332 AVSS 0.089409f
C7638 AVDD.t1199 AVSS 0.089409f
C7639 AVDD.n460 AVSS 0.342362f
C7640 AVDD.t569 AVSS 0.089409f
C7641 AVDD.t150 AVSS 0.089409f
C7642 AVDD.n461 AVSS 0.261503f
C7643 AVDD.t570 AVSS 0.045717f
C7644 AVDD.t1004 AVSS 0.045717f
C7645 AVDD.n462 AVSS 0.284944f
C7646 AVDD.t1003 AVSS 0.089409f
C7647 AVDD.n463 AVSS 0.225482f
C7648 AVDD.t635 AVSS 0.089409f
C7649 AVDD.n464 AVSS 0.225482f
C7650 AVDD.t636 AVSS 0.045717f
C7651 AVDD.n465 AVSS 0.376621f
C7652 AVDD.t1256 AVSS 0.045717f
C7653 AVDD.t100 AVSS 0.089409f
C7654 AVDD.n466 AVSS 0.225482f
C7655 AVDD.t1255 AVSS 0.089409f
C7656 AVDD.n467 AVSS 0.225482f
C7657 AVDD.n468 AVSS 0.376621f
C7658 AVDD.n469 AVSS 0.68361f
C7659 AVDD.n470 AVSS 0.236716f
C7660 AVDD.t151 AVSS 0.045717f
C7661 AVDD.n471 AVSS 0.320025f
C7662 AVDD.n472 AVSS 0.320025f
C7663 AVDD.t333 AVSS 0.033572f
C7664 AVDD.n473 AVSS 0.021426f
C7665 AVDD.n474 AVSS 0.278352f
C7666 AVDD.n475 AVSS 0.021426f
C7667 AVDD.t940 AVSS 0.021426f
C7668 AVDD.n476 AVSS 0.021426f
C7669 AVDD.n477 AVSS 0.278352f
C7670 AVDD.n478 AVSS 0.021426f
C7671 AVDD.t1022 AVSS 0.021426f
C7672 AVDD.n479 AVSS 0.021426f
C7673 AVDD.n480 AVSS 0.278352f
C7674 AVDD.n481 AVSS 0.021426f
C7675 AVDD.t348 AVSS 0.033572f
C7676 AVDD.n482 AVSS 0.292092f
C7677 AVDD.n483 AVSS 0.292092f
C7678 AVDD.t382 AVSS 0.033572f
C7679 AVDD.n484 AVSS 0.021426f
C7680 AVDD.n485 AVSS 0.26267f
C7681 AVDD.n486 AVSS 0.021426f
C7682 AVDD.t364 AVSS 0.021426f
C7683 AVDD.n487 AVSS 0.021426f
C7684 AVDD.n488 AVSS 0.278352f
C7685 AVDD.n489 AVSS 0.021426f
C7686 AVDD.t970 AVSS 0.033572f
C7687 AVDD.n490 AVSS 0.292092f
C7688 AVDD.n491 AVSS 0.292092f
C7689 AVDD.t1078 AVSS 0.033572f
C7690 AVDD.n492 AVSS 0.021426f
C7691 AVDD.n493 AVSS 0.278352f
C7692 AVDD.n494 AVSS 0.021426f
C7693 AVDD.t280 AVSS 0.021426f
C7694 AVDD.n495 AVSS 0.021426f
C7695 AVDD.n496 AVSS 0.278352f
C7696 AVDD.n497 AVSS 0.021426f
C7697 AVDD.t292 AVSS 0.021426f
C7698 AVDD.n498 AVSS 0.021426f
C7699 AVDD.n499 AVSS 0.278352f
C7700 AVDD.n500 AVSS 0.021426f
C7701 AVDD.t736 AVSS 0.033572f
C7702 AVDD.n501 AVSS 0.301403f
C7703 AVDD.n502 AVSS 0.763137f
C7704 AVDD.t1002 AVSS 0.045717f
C7705 AVDD.t582 AVSS 0.045717f
C7706 AVDD.n503 AVSS 0.446192f
C7707 AVDD.t581 AVSS 0.089409f
C7708 AVDD.t1001 AVSS 0.089409f
C7709 AVDD.n504 AVSS 0.787444f
C7710 AVDD.t420 AVSS 0.045717f
C7711 AVDD.t1258 AVSS 0.045717f
C7712 AVDD.n505 AVSS 0.764636f
C7713 AVDD.t1257 AVSS 0.089409f
C7714 AVDD.t419 AVSS 0.089409f
C7715 AVDD.n506 AVSS 0.445699f
C7716 AVDD.t108 AVSS 0.089409f
C7717 AVDD.t544 AVSS 0.089409f
C7718 AVDD.n507 AVSS 0.445699f
C7719 AVDD.t545 AVSS 0.045717f
C7720 AVDD.t109 AVSS 0.045717f
C7721 AVDD.n508 AVSS 0.537731f
C7722 AVDD.n509 AVSS 0.378581f
C7723 AVDD.n510 AVSS 0.712338f
C7724 AVDD.t529 AVSS 0.045717f
C7725 AVDD.t80 AVSS 0.045717f
C7726 AVDD.n511 AVSS 0.587661f
C7727 AVDD.t78 AVSS 0.089409f
C7728 AVDD.t528 AVSS 0.089409f
C7729 AVDD.n512 AVSS 0.445699f
C7730 AVDD.t213 AVSS 0.089409f
C7731 AVDD.t633 AVSS 0.089409f
C7732 AVDD.n513 AVSS 0.445699f
C7733 AVDD.t634 AVSS 0.045717f
C7734 AVDD.t214 AVSS 0.045717f
C7735 AVDD.n514 AVSS 0.764636f
C7736 AVDD.t989 AVSS 0.089409f
C7737 AVDD.t126 AVSS 0.089409f
C7738 AVDD.n515 AVSS 0.787444f
C7739 AVDD.t127 AVSS 0.045717f
C7740 AVDD.t990 AVSS 0.045717f
C7741 AVDD.n516 AVSS 0.23704f
C7742 AVDD.n517 AVSS 0.608466f
C7743 AVDD.n518 AVSS 0.153168f
C7744 AVDD.t274 AVSS 0.089409f
C7745 AVDD.n519 AVSS 0.173626f
C7746 AVDD.n520 AVSS 0.141621f
C7747 AVDD.n521 AVSS 0.021426f
C7748 AVDD.t689 AVSS 0.021426f
C7749 AVDD.n522 AVSS 0.021426f
C7750 AVDD.n523 AVSS 0.141621f
C7751 AVDD.t1061 AVSS 0.089409f
C7752 AVDD.n524 AVSS 0.173626f
C7753 AVDD.n525 AVSS 0.141621f
C7754 AVDD.n526 AVSS 0.021426f
C7755 AVDD.t218 AVSS 0.033572f
C7756 AVDD.n527 AVSS 0.148431f
C7757 AVDD.n528 AVSS 0.148431f
C7758 AVDD.t491 AVSS 0.033572f
C7759 AVDD.n529 AVSS 0.021426f
C7760 AVDD.n530 AVSS 0.141621f
C7761 AVDD.t791 AVSS 0.089409f
C7762 AVDD.n531 AVSS 0.110794f
C7763 AVDD.n532 AVSS 0.07081f
C7764 AVDD.n533 AVSS 0.133642f
C7765 AVDD.n534 AVSS 0.021426f
C7766 AVDD.t1190 AVSS 0.033572f
C7767 AVDD.n535 AVSS 0.148431f
C7768 AVDD.n536 AVSS 0.148431f
C7769 AVDD.t1159 AVSS 0.089409f
C7770 AVDD.n537 AVSS 0.173626f
C7771 AVDD.n538 AVSS 0.141621f
C7772 AVDD.n539 AVSS 0.021426f
C7773 AVDD.t134 AVSS 0.021426f
C7774 AVDD.n540 AVSS 0.021426f
C7775 AVDD.n541 AVSS 0.141621f
C7776 AVDD.t445 AVSS 0.089409f
C7777 AVDD.n542 AVSS 0.173626f
C7778 AVDD.n543 AVSS 0.141621f
C7779 AVDD.n544 AVSS 0.021426f
C7780 AVDD.t750 AVSS 0.033572f
C7781 AVDD.n545 AVSS 0.197553f
C7782 AVDD.n546 AVSS 0.38292f
C7783 AVDD.t979 AVSS 0.089409f
C7784 AVDD.n547 AVSS 0.398711f
C7785 AVDD.n548 AVSS 0.387307f
C7786 AVDD.t202 AVSS 0.089409f
C7787 AVDD.n549 AVSS 0.225482f
C7788 AVDD.t66 AVSS 0.089409f
C7789 AVDD.n550 AVSS 0.225482f
C7790 AVDD.n551 AVSS 0.218015f
C7791 AVDD.n552 AVSS 0.196027f
C7792 AVDD.n553 AVSS 0.24747f
C7793 AVDD.n554 AVSS 0.375467f
C7794 AVDD.t347 AVSS 12.609f
C7795 AVDD.t122 AVSS 10.1876f
C7796 AVDD.t19 AVSS 10.1876f
C7797 AVDD.t44 AVSS 13.1202f
C7798 AVDD.t67 AVSS 12.2951f
C7799 AVDD.n555 AVSS 6.02649f
C7800 AVDD.n556 AVSS 0.375467f
C7801 AVDD.n557 AVSS 0.180541f
C7802 AVDD.n558 AVSS 0.27229f
C7803 AVDD.t997 AVSS 0.089409f
C7804 AVDD.n559 AVSS 0.225482f
C7805 AVDD.t1093 AVSS 0.089409f
C7806 AVDD.n560 AVSS 0.225482f
C7807 AVDD.n561 AVSS 0.376621f
C7808 AVDD.n562 AVSS 0.789554f
C7809 AVDD.n563 AVSS 0.401227f
C7810 AVDD.t592 AVSS 0.045717f
C7811 AVDD.n564 AVSS 0.547954f
C7812 AVDD.n565 AVSS 0.547954f
C7813 AVDD.t829 AVSS 0.033572f
C7814 AVDD.n566 AVSS 0.021426f
C7815 AVDD.n567 AVSS 0.49024f
C7816 AVDD.n568 AVSS 0.021426f
C7817 AVDD.t768 AVSS 0.021426f
C7818 AVDD.n569 AVSS 0.021426f
C7819 AVDD.n570 AVSS 0.49024f
C7820 AVDD.n571 AVSS 0.021426f
C7821 AVDD.t1274 AVSS 0.021426f
C7822 AVDD.n572 AVSS 0.021426f
C7823 AVDD.n573 AVSS 0.49024f
C7824 AVDD.n574 AVSS 0.021426f
C7825 AVDD.t1224 AVSS 0.033572f
C7826 AVDD.n575 AVSS 0.498758f
C7827 AVDD.n576 AVSS 0.498758f
C7828 AVDD.t531 AVSS 0.033572f
C7829 AVDD.n577 AVSS 0.021426f
C7830 AVDD.n578 AVSS 0.462621f
C7831 AVDD.n579 AVSS 0.021426f
C7832 AVDD.t914 AVSS 0.021426f
C7833 AVDD.n580 AVSS 0.021426f
C7834 AVDD.n581 AVSS 0.49024f
C7835 AVDD.n582 AVSS 0.021426f
C7836 AVDD.t859 AVSS 0.033572f
C7837 AVDD.n583 AVSS 0.498758f
C7838 AVDD.n584 AVSS 0.498758f
C7839 AVDD.t468 AVSS 0.033572f
C7840 AVDD.n585 AVSS 0.021426f
C7841 AVDD.n586 AVSS 0.49024f
C7842 AVDD.n587 AVSS 0.021426f
C7843 AVDD.t857 AVSS 0.021426f
C7844 AVDD.n588 AVSS 0.021426f
C7845 AVDD.n589 AVSS 0.49024f
C7846 AVDD.n590 AVSS 0.021426f
C7847 AVDD.t788 AVSS 0.021426f
C7848 AVDD.n591 AVSS 0.021426f
C7849 AVDD.n592 AVSS 0.49024f
C7850 AVDD.n593 AVSS 0.021426f
C7851 AVDD.t1148 AVSS 0.033572f
C7852 AVDD.n594 AVSS 0.547954f
C7853 AVDD.n595 AVSS 0.547954f
C7854 AVDD.t408 AVSS 0.045717f
C7855 AVDD.n596 AVSS 0.493579f
C7856 AVDD.n597 AVSS 1.52977f
C7857 AVDD.n598 AVSS 0.493579f
C7858 AVDD.t968 AVSS 0.045717f
C7859 AVDD.n599 AVSS 0.547954f
C7860 AVDD.n600 AVSS 0.547954f
C7861 AVDD.t250 AVSS 0.033572f
C7862 AVDD.n601 AVSS 0.021426f
C7863 AVDD.n602 AVSS 0.49024f
C7864 AVDD.n603 AVSS 0.021426f
C7865 AVDD.t165 AVSS 0.021426f
C7866 AVDD.n604 AVSS 0.021426f
C7867 AVDD.n605 AVSS 0.49024f
C7868 AVDD.n606 AVSS 0.021426f
C7869 AVDD.t541 AVSS 0.021426f
C7870 AVDD.n607 AVSS 0.021426f
C7871 AVDD.n608 AVSS 0.49024f
C7872 AVDD.n609 AVSS 0.021426f
C7873 AVDD.t462 AVSS 0.033572f
C7874 AVDD.n610 AVSS 0.498758f
C7875 AVDD.t236 AVSS 0.021426f
C7876 AVDD.n611 AVSS 0.021426f
C7877 AVDD.t1152 AVSS 0.033572f
C7878 AVDD.t1151 AVSS 0.089409f
C7879 AVDD.t1145 AVSS 0.089409f
C7880 AVDD.n612 AVSS 0.55425f
C7881 AVDD.n613 AVSS 0.498758f
C7882 AVDD.t1146 AVSS 0.033572f
C7883 AVDD.n614 AVSS 0.021426f
C7884 AVDD.t231 AVSS 0.021426f
C7885 AVDD.t161 AVSS 0.033572f
C7886 AVDD.t770 AVSS 0.033572f
C7887 AVDD.t769 AVSS 0.089409f
C7888 AVDD.t761 AVSS 0.089409f
C7889 AVDD.n615 AVSS 0.55425f
C7890 AVDD.t1110 AVSS 0.021426f
C7891 AVDD.n616 AVSS 0.021426f
C7892 AVDD.t1117 AVSS 0.089409f
C7893 AVDD.t1118 AVSS 0.021426f
C7894 AVDD.n617 AVSS 0.021426f
C7895 AVDD.t1047 AVSS 0.089409f
C7896 AVDD.t1039 AVSS 0.089409f
C7897 AVDD.n618 AVSS 0.55425f
C7898 AVDD.t454 AVSS 0.033572f
C7899 AVDD.t1048 AVSS 0.021426f
C7900 AVDD.n619 AVSS 0.021426f
C7901 AVDD.t463 AVSS 0.089409f
C7902 AVDD.t464 AVSS 0.033572f
C7903 AVDD.t1216 AVSS 0.033572f
C7904 AVDD.t1215 AVSS 0.089409f
C7905 AVDD.t1209 AVSS 0.089409f
C7906 AVDD.n620 AVSS 0.55425f
C7907 AVDD.t1126 AVSS 0.021426f
C7908 AVDD.n621 AVSS 0.021426f
C7909 AVDD.t1133 AVSS 0.089409f
C7910 AVDD.t1134 AVSS 0.021426f
C7911 AVDD.n622 AVSS 0.021426f
C7912 AVDD.t1045 AVSS 0.089409f
C7913 AVDD.t1035 AVSS 0.089409f
C7914 AVDD.n623 AVSS 0.55425f
C7915 AVDD.t594 AVSS 0.033572f
C7916 AVDD.t1046 AVSS 0.021426f
C7917 AVDD.n624 AVSS 0.021426f
C7918 AVDD.t599 AVSS 0.089409f
C7919 AVDD.t600 AVSS 0.033572f
C7920 AVDD.t11 AVSS 0.033572f
C7921 AVDD.t10 AVSS 0.089409f
C7922 AVDD.t4 AVSS 0.089409f
C7923 AVDD.n625 AVSS 0.55425f
C7924 AVDD.t99 AVSS 0.021426f
C7925 AVDD.n626 AVSS 0.021426f
C7926 AVDD.t106 AVSS 0.089409f
C7927 AVDD.t107 AVSS 0.021426f
C7928 AVDD.n627 AVSS 0.021426f
C7929 AVDD.t1019 AVSS 0.089409f
C7930 AVDD.t1015 AVSS 0.089409f
C7931 AVDD.n628 AVSS 0.55425f
C7932 AVDD.t1020 AVSS 0.033572f
C7933 AVDD.t430 AVSS 0.033572f
C7934 AVDD.t429 AVSS 0.089409f
C7935 AVDD.t425 AVSS 0.089409f
C7936 AVDD.n629 AVSS 0.55425f
C7937 AVDD.t495 AVSS 0.021426f
C7938 AVDD.n630 AVSS 0.021426f
C7939 AVDD.t502 AVSS 0.089409f
C7940 AVDD.t503 AVSS 0.021426f
C7941 AVDD.n631 AVSS 0.021426f
C7942 AVDD.t1081 AVSS 0.089409f
C7943 AVDD.t1067 AVSS 0.089409f
C7944 AVDD.n632 AVSS 0.55425f
C7945 AVDD.t1158 AVSS 0.033572f
C7946 AVDD.t1082 AVSS 0.021426f
C7947 AVDD.n633 AVSS 0.021426f
C7948 AVDD.t1165 AVSS 0.089409f
C7949 AVDD.t1166 AVSS 0.033572f
C7950 AVDD.t942 AVSS 0.045717f
C7951 AVDD.t941 AVSS 0.089409f
C7952 AVDD.t937 AVSS 0.089409f
C7953 AVDD.n634 AVSS 0.55425f
C7954 AVDD.t566 AVSS 0.045717f
C7955 AVDD.t144 AVSS 0.045717f
C7956 AVDD.n635 AVSS 0.743554f
C7957 AVDD.t25 AVSS 0.045717f
C7958 AVDD.t24 AVSS 0.089409f
C7959 AVDD.t7 AVSS 0.089409f
C7960 AVDD.n636 AVSS 0.55425f
C7961 AVDD.t1104 AVSS 0.033572f
C7962 AVDD.t1103 AVSS 0.089409f
C7963 AVDD.t1097 AVSS 0.089409f
C7964 AVDD.n637 AVSS 0.55425f
C7965 AVDD.t748 AVSS 0.021426f
C7966 AVDD.n638 AVSS 0.021426f
C7967 AVDD.t755 AVSS 0.089409f
C7968 AVDD.t756 AVSS 0.021426f
C7969 AVDD.n639 AVSS 0.021426f
C7970 AVDD.t484 AVSS 0.089409f
C7971 AVDD.t471 AVSS 0.089409f
C7972 AVDD.n640 AVSS 0.55425f
C7973 AVDD.t91 AVSS 0.033572f
C7974 AVDD.t485 AVSS 0.021426f
C7975 AVDD.n641 AVSS 0.021426f
C7976 AVDD.t102 AVSS 0.089409f
C7977 AVDD.t103 AVSS 0.033572f
C7978 AVDD.t509 AVSS 0.033572f
C7979 AVDD.t508 AVSS 0.089409f
C7980 AVDD.t500 AVSS 0.089409f
C7981 AVDD.n642 AVSS 0.55425f
C7982 AVDD.t906 AVSS 0.021426f
C7983 AVDD.n643 AVSS 0.021426f
C7984 AVDD.n644 AVSS 0.374271f
C7985 AVDD.t911 AVSS 0.089409f
C7986 AVDD.t912 AVSS 0.021426f
C7987 AVDD.n645 AVSS 0.021426f
C7988 AVDD.t532 AVSS 0.089409f
C7989 AVDD.t526 AVSS 0.089409f
C7990 AVDD.n646 AVSS 0.55425f
C7991 AVDD.t533 AVSS 0.033572f
C7992 AVDD.t910 AVSS 0.033572f
C7993 AVDD.t909 AVSS 0.089409f
C7994 AVDD.t903 AVSS 0.089409f
C7995 AVDD.n647 AVSS 0.55425f
C7996 AVDD.t966 AVSS 0.021426f
C7997 AVDD.n648 AVSS 0.021426f
C7998 AVDD.t971 AVSS 0.089409f
C7999 AVDD.t972 AVSS 0.021426f
C8000 AVDD.n649 AVSS 0.021426f
C8001 AVDD.t288 AVSS 0.089409f
C8002 AVDD.t284 AVSS 0.089409f
C8003 AVDD.n650 AVSS 0.55425f
C8004 AVDD.t665 AVSS 0.033572f
C8005 AVDD.t289 AVSS 0.021426f
C8006 AVDD.n651 AVSS 0.021426f
C8007 AVDD.t672 AVSS 0.089409f
C8008 AVDD.t673 AVSS 0.033572f
C8009 AVDD.t117 AVSS 0.045717f
C8010 AVDD.t116 AVSS 0.089409f
C8011 AVDD.t104 AVSS 0.089409f
C8012 AVDD.n652 AVSS 0.402345f
C8013 AVDD.t833 AVSS 0.045717f
C8014 AVDD.n653 AVSS 0.367741f
C8015 AVDD.t626 AVSS 0.045717f
C8016 AVDD.t515 AVSS 0.045717f
C8017 AVDD.t521 AVSS 0.045717f
C8018 AVDD.n654 AVSS 0.29069f
C8019 AVDD.n655 AVSS 0.378609f
C8020 AVDD.t62 AVSS 12.2951f
C8021 AVDD.n656 AVSS 0.378581f
C8022 AVDD.n657 AVSS 0.374271f
C8023 AVDD.n658 AVSS 0.378609f
C8024 AVDD.t414 AVSS 0.045717f
C8025 AVDD.n659 AVSS 0.266012f
C8026 AVDD.t406 AVSS 0.045717f
C8027 AVDD.t517 AVSS 0.045717f
C8028 AVDD.t1262 AVSS 0.045717f
C8029 AVDD.t739 AVSS 0.089409f
C8030 AVDD.n660 AVSS 0.173626f
C8031 AVDD.t790 AVSS 0.021426f
C8032 AVDD.n661 AVSS 0.342168f
C8033 AVDD.t922 AVSS 0.033572f
C8034 AVDD.t655 AVSS 0.045717f
C8035 AVDD.n662 AVSS 0.342168f
C8036 AVDD.t984 AVSS 0.045717f
C8037 AVDD.n663 AVSS 0.206516f
C8038 AVDD.n664 AVSS 0.464086f
C8039 AVDD.t946 AVSS 0.045717f
C8040 AVDD.t132 AVSS 0.045717f
C8041 AVDD.t678 AVSS 0.089409f
C8042 AVDD.n665 AVSS 0.207359f
C8043 AVDD.n666 AVSS 0.006326f
C8044 AVDD.t1646 AVSS 0.010713f
C8045 AVDD.t1481 AVSS 0.010713f
C8046 AVDD.n667 AVSS 0.024349f
C8047 AVDD.n668 AVSS 0.020751f
C8048 AVDD.n669 AVSS 0.006326f
C8049 AVDD.t1380 AVSS 0.010713f
C8050 AVDD.t1412 AVSS 0.010713f
C8051 AVDD.n670 AVSS 0.024349f
C8052 AVDD.n671 AVSS 0.020751f
C8053 AVDD.n672 AVSS 0.006326f
C8054 AVDD.t1663 AVSS 0.025767f
C8055 AVDD.n673 AVSS 0.031066f
C8056 AVDD.n674 AVSS 0.006326f
C8057 AVDD.t1471 AVSS 0.010713f
C8058 AVDD.t1444 AVSS 0.010713f
C8059 AVDD.n675 AVSS 0.024349f
C8060 AVDD.n676 AVSS 0.020751f
C8061 AVDD.n677 AVSS 0.006326f
C8062 AVDD.t1287 AVSS 0.010713f
C8063 AVDD.t1595 AVSS 0.010713f
C8064 AVDD.n678 AVSS 0.024349f
C8065 AVDD.n679 AVSS 0.020751f
C8066 AVDD.n680 AVSS 0.006326f
C8067 AVDD.t1407 AVSS 0.010713f
C8068 AVDD.t1298 AVSS 0.010713f
C8069 AVDD.n681 AVSS 0.024349f
C8070 AVDD.n682 AVSS 0.020751f
C8071 AVDD.t983 AVSS 0.089409f
C8072 AVDD.n683 AVSS 0.218463f
C8073 AVDD.t180 AVSS 0.089409f
C8074 AVDD.n684 AVSS 0.218463f
C8075 AVDD.t182 AVSS 0.045717f
C8076 AVDD.n685 AVSS 0.194592f
C8077 AVDD.t724 AVSS 0.045717f
C8078 AVDD.n686 AVSS 0.147702f
C8079 AVDD.n687 AVSS 0.006326f
C8080 AVDD.n688 AVSS 0.006326f
C8081 AVDD.n689 AVSS 0.006326f
C8082 AVDD.n690 AVSS 0.006326f
C8083 AVDD.n691 AVSS 0.006326f
C8084 AVDD.n692 AVSS 0.006326f
C8085 AVDD.t679 AVSS 0.045717f
C8086 AVDD.n693 AVSS 0.211203f
C8087 AVDD.t1080 AVSS 0.045717f
C8088 AVDD.n694 AVSS 0.31086f
C8089 AVDD.n695 AVSS 0.292136f
C8090 AVDD.t1121 AVSS 0.089409f
C8091 AVDD.n696 AVSS 0.363872f
C8092 AVDD.t657 AVSS 0.021426f
C8093 AVDD.t511 AVSS 0.033572f
C8094 AVDD.t64 AVSS 0.089409f
C8095 AVDD.n697 AVSS 0.363872f
C8096 AVDD.n698 AVSS 0.331867f
C8097 AVDD.n699 AVSS 0.336325f
C8098 AVDD.t367 AVSS 0.021426f
C8099 AVDD.t272 AVSS 0.089409f
C8100 AVDD.n700 AVSS 0.363872f
C8101 AVDD.t365 AVSS 0.089409f
C8102 AVDD.n701 AVSS 0.326478f
C8103 AVDD.t1251 AVSS 0.089409f
C8104 AVDD.n702 AVSS 0.363872f
C8105 AVDD.n703 AVSS 0.331651f
C8106 AVDD.t273 AVSS 0.033572f
C8107 AVDD.t641 AVSS 0.033572f
C8108 AVDD.n704 AVSS 0.326024f
C8109 AVDD.t215 AVSS 0.089409f
C8110 AVDD.n705 AVSS 0.075241f
C8111 AVDD.n706 AVSS 0.331867f
C8112 AVDD.n707 AVSS 0.342167f
C8113 AVDD.n708 AVSS 0.021426f
C8114 AVDD.t744 AVSS 0.021426f
C8115 AVDD.t1203 AVSS 0.089409f
C8116 AVDD.n709 AVSS 0.347512f
C8117 AVDD.n710 AVSS 0.342167f
C8118 AVDD.t921 AVSS 0.089409f
C8119 AVDD.n711 AVSS 0.41412f
C8120 AVDD.n712 AVSS 0.342167f
C8121 AVDD.t1204 AVSS 0.033572f
C8122 AVDD.n713 AVSS 0.021426f
C8123 AVDD.n714 AVSS 0.331867f
C8124 AVDD.t640 AVSS 0.089409f
C8125 AVDD.n715 AVSS 0.363872f
C8126 AVDD.t743 AVSS 0.089409f
C8127 AVDD.n716 AVSS 0.363872f
C8128 AVDD.n717 AVSS 0.331867f
C8129 AVDD.n718 AVSS 0.021426f
C8130 AVDD.t216 AVSS 0.021426f
C8131 AVDD.n719 AVSS 0.021426f
C8132 AVDD.n720 AVSS 0.331867f
C8133 AVDD.n721 AVSS 0.331867f
C8134 AVDD.n722 AVSS 0.021426f
C8135 AVDD.t1252 AVSS 0.033572f
C8136 AVDD.n723 AVSS 0.336325f
C8137 AVDD.t228 AVSS 0.089409f
C8138 AVDD.n724 AVSS 0.347512f
C8139 AVDD.t656 AVSS 0.089409f
C8140 AVDD.n725 AVSS 0.363872f
C8141 AVDD.t26 AVSS 0.089409f
C8142 AVDD.n726 AVSS 0.363872f
C8143 AVDD.t686 AVSS 0.089409f
C8144 AVDD.n727 AVSS 0.41412f
C8145 AVDD.t902 AVSS 0.021426f
C8146 AVDD.t1249 AVSS 0.089409f
C8147 AVDD.n728 AVSS 0.363872f
C8148 AVDD.t1088 AVSS 0.033572f
C8149 AVDD.t1087 AVSS 0.089409f
C8150 AVDD.t708 AVSS 0.089409f
C8151 AVDD.n729 AVSS 0.342362f
C8152 AVDD.t1124 AVSS 0.021426f
C8153 AVDD.n730 AVSS 0.021426f
C8154 AVDD.t254 AVSS 0.089409f
C8155 AVDD.t256 AVSS 0.021426f
C8156 AVDD.n731 AVSS 0.021426f
C8157 AVDD.t955 AVSS 0.089409f
C8158 AVDD.t561 AVSS 0.089409f
C8159 AVDD.n732 AVSS 0.342362f
C8160 AVDD.t986 AVSS 0.033572f
C8161 AVDD.t956 AVSS 0.021426f
C8162 AVDD.n733 AVSS 0.021426f
C8163 AVDD.t81 AVSS 0.089409f
C8164 AVDD.t83 AVSS 0.033572f
C8165 AVDD.t1138 AVSS 0.033572f
C8166 AVDD.t1137 AVSS 0.089409f
C8167 AVDD.t733 AVSS 0.089409f
C8168 AVDD.n734 AVSS 0.342362f
C8169 AVDD.t697 AVSS 0.021426f
C8170 AVDD.n735 AVSS 0.021426f
C8171 AVDD.t1071 AVSS 0.089409f
C8172 AVDD.t1072 AVSS 0.021426f
C8173 AVDD.n736 AVSS 0.021426f
C8174 AVDD.t232 AVSS 0.089409f
C8175 AVDD.t1101 AVSS 0.089409f
C8176 AVDD.n737 AVSS 0.342362f
C8177 AVDD.t234 AVSS 0.033572f
C8178 AVDD.t507 AVSS 0.033572f
C8179 AVDD.t506 AVSS 0.089409f
C8180 AVDD.t92 AVSS 0.089409f
C8181 AVDD.n738 AVSS 0.342362f
C8182 AVDD.t379 AVSS 0.021426f
C8183 AVDD.n739 AVSS 0.021426f
C8184 AVDD.t801 AVSS 0.089409f
C8185 AVDD.t802 AVSS 0.021426f
C8186 AVDD.n740 AVSS 0.021426f
C8187 AVDD.t361 AVSS 0.089409f
C8188 AVDD.t1231 AVSS 0.089409f
C8189 AVDD.n741 AVSS 0.342362f
C8190 AVDD.t1198 AVSS 0.033572f
C8191 AVDD.t362 AVSS 0.021426f
C8192 AVDD.n742 AVSS 0.021426f
C8193 AVDD.t325 AVSS 0.089409f
C8194 AVDD.t326 AVSS 0.033572f
C8195 AVDD.t896 AVSS 0.045717f
C8196 AVDD.t895 AVSS 0.089409f
C8197 AVDD.t477 AVSS 0.089409f
C8198 AVDD.n743 AVSS 0.256112f
C8199 AVDD.t313 AVSS 0.045717f
C8200 AVDD.t413 AVSS 0.089409f
C8201 AVDD.n744 AVSS 0.220656f
C8202 AVDD.t312 AVSS 0.089409f
C8203 AVDD.n745 AVSS 0.220656f
C8204 AVDD.n746 AVSS 0.367741f
C8205 AVDD.t520 AVSS 0.089409f
C8206 AVDD.n747 AVSS 0.220656f
C8207 AVDD.t1195 AVSS 0.089409f
C8208 AVDD.n748 AVSS 0.220656f
C8209 AVDD.t1196 AVSS 0.045717f
C8210 AVDD.n749 AVSS 0.367741f
C8211 AVDD.n750 AVSS 0.670031f
C8212 AVDD.n751 AVSS 0.3558f
C8213 AVDD.t478 AVSS 0.045717f
C8214 AVDD.n752 AVSS 0.320025f
C8215 AVDD.n753 AVSS 0.320025f
C8216 AVDD.t1197 AVSS 0.089409f
C8217 AVDD.n754 AVSS 0.342362f
C8218 AVDD.n755 AVSS 0.278352f
C8219 AVDD.n756 AVSS 0.021426f
C8220 AVDD.t1232 AVSS 0.021426f
C8221 AVDD.n757 AVSS 0.021426f
C8222 AVDD.n758 AVSS 0.278352f
C8223 AVDD.t377 AVSS 0.089409f
C8224 AVDD.n759 AVSS 0.342362f
C8225 AVDD.n760 AVSS 0.278352f
C8226 AVDD.n761 AVSS 0.021426f
C8227 AVDD.t94 AVSS 0.033572f
C8228 AVDD.n762 AVSS 0.292092f
C8229 AVDD.n763 AVSS 0.292092f
C8230 AVDD.t1102 AVSS 0.033572f
C8231 AVDD.n764 AVSS 0.021426f
C8232 AVDD.n765 AVSS 0.278352f
C8233 AVDD.t696 AVSS 0.089409f
C8234 AVDD.n766 AVSS 0.218868f
C8235 AVDD.n767 AVSS 0.139176f
C8236 AVDD.n768 AVSS 0.26267f
C8237 AVDD.n769 AVSS 0.021426f
C8238 AVDD.t734 AVSS 0.033572f
C8239 AVDD.n770 AVSS 0.292092f
C8240 AVDD.n771 AVSS 0.292092f
C8241 AVDD.t985 AVSS 0.089409f
C8242 AVDD.n772 AVSS 0.342362f
C8243 AVDD.n773 AVSS 0.278352f
C8244 AVDD.n774 AVSS 0.021426f
C8245 AVDD.t562 AVSS 0.021426f
C8246 AVDD.n775 AVSS 0.021426f
C8247 AVDD.n776 AVSS 0.278352f
C8248 AVDD.t1123 AVSS 0.089409f
C8249 AVDD.n777 AVSS 0.342362f
C8250 AVDD.n778 AVSS 0.278352f
C8251 AVDD.n779 AVSS 0.021426f
C8252 AVDD.t709 AVSS 0.033572f
C8253 AVDD.n780 AVSS 0.301403f
C8254 AVDD.t745 AVSS 0.089409f
C8255 AVDD.t334 AVSS 0.089409f
C8256 AVDD.n781 AVSS 0.342362f
C8257 AVDD.t746 AVSS 0.033572f
C8258 AVDD.t31 AVSS 0.021426f
C8259 AVDD.t443 AVSS 0.089409f
C8260 AVDD.t29 AVSS 0.089409f
C8261 AVDD.n782 AVSS 0.342362f
C8262 AVDD.t892 AVSS 0.021426f
C8263 AVDD.t891 AVSS 0.089409f
C8264 AVDD.t469 AVSS 0.089409f
C8265 AVDD.n783 AVSS 0.342362f
C8266 AVDD.t196 AVSS 0.033572f
C8267 AVDD.t601 AVSS 0.089409f
C8268 AVDD.t195 AVSS 0.089409f
C8269 AVDD.n784 AVSS 0.342362f
C8270 AVDD.t646 AVSS 0.089409f
C8271 AVDD.t251 AVSS 0.089409f
C8272 AVDD.n785 AVSS 0.342362f
C8273 AVDD.t647 AVSS 0.033572f
C8274 AVDD.t1086 AVSS 0.021426f
C8275 AVDD.t219 AVSS 0.089409f
C8276 AVDD.t1085 AVSS 0.089409f
C8277 AVDD.n786 AVSS 0.218868f
C8278 AVDD.t1212 AVSS 0.033572f
C8279 AVDD.t1211 AVSS 0.089409f
C8280 AVDD.t834 AVSS 0.089409f
C8281 AVDD.n787 AVSS 0.342362f
C8282 AVDD.n788 AVSS 0.139176f
C8283 AVDD.t1053 AVSS 0.089409f
C8284 AVDD.t662 AVSS 0.089409f
C8285 AVDD.n789 AVSS 0.342362f
C8286 AVDD.t1054 AVSS 0.033572f
C8287 AVDD.t645 AVSS 0.021426f
C8288 AVDD.t1031 AVSS 0.089409f
C8289 AVDD.t644 AVSS 0.089409f
C8290 AVDD.n790 AVSS 0.342362f
C8291 AVDD.t142 AVSS 0.021426f
C8292 AVDD.t140 AVSS 0.089409f
C8293 AVDD.t1025 AVSS 0.089409f
C8294 AVDD.n791 AVSS 0.342362f
C8295 AVDD.t295 AVSS 0.033572f
C8296 AVDD.t682 AVSS 0.089409f
C8297 AVDD.t293 AVSS 0.089409f
C8298 AVDD.n792 AVSS 0.342362f
C8299 AVDD.t683 AVSS 0.033572f
C8300 AVDD.n793 AVSS 0.021426f
C8301 AVDD.n794 AVSS 0.278352f
C8302 AVDD.n795 AVSS 0.021426f
C8303 AVDD.t1026 AVSS 0.021426f
C8304 AVDD.n796 AVSS 0.021426f
C8305 AVDD.n797 AVSS 0.278352f
C8306 AVDD.n798 AVSS 0.021426f
C8307 AVDD.t1032 AVSS 0.021426f
C8308 AVDD.n799 AVSS 0.021426f
C8309 AVDD.n800 AVSS 0.278352f
C8310 AVDD.n801 AVSS 0.021426f
C8311 AVDD.t663 AVSS 0.033572f
C8312 AVDD.n802 AVSS 0.292092f
C8313 AVDD.n803 AVSS 0.292092f
C8314 AVDD.t835 AVSS 0.033572f
C8315 AVDD.n804 AVSS 0.021426f
C8316 AVDD.n805 AVSS 0.26267f
C8317 AVDD.n806 AVSS 0.021426f
C8318 AVDD.t220 AVSS 0.021426f
C8319 AVDD.n807 AVSS 0.021426f
C8320 AVDD.n808 AVSS 0.278352f
C8321 AVDD.n809 AVSS 0.021426f
C8322 AVDD.t253 AVSS 0.033572f
C8323 AVDD.n810 AVSS 0.292092f
C8324 AVDD.n811 AVSS 0.292092f
C8325 AVDD.t602 AVSS 0.033572f
C8326 AVDD.n812 AVSS 0.021426f
C8327 AVDD.n813 AVSS 0.278352f
C8328 AVDD.n814 AVSS 0.021426f
C8329 AVDD.t470 AVSS 0.021426f
C8330 AVDD.n815 AVSS 0.021426f
C8331 AVDD.n816 AVSS 0.278352f
C8332 AVDD.n817 AVSS 0.021426f
C8333 AVDD.t444 AVSS 0.021426f
C8334 AVDD.n818 AVSS 0.021426f
C8335 AVDD.n819 AVSS 0.278352f
C8336 AVDD.n820 AVSS 0.021426f
C8337 AVDD.t336 AVSS 0.033572f
C8338 AVDD.n821 AVSS 0.301403f
C8339 AVDD.t143 AVSS 0.089409f
C8340 AVDD.t565 AVSS 0.089409f
C8341 AVDD.n822 AVSS 0.445699f
C8342 AVDD.t15 AVSS 0.089409f
C8343 AVDD.t437 AVSS 0.089409f
C8344 AVDD.n823 AVSS 0.445699f
C8345 AVDD.t438 AVSS 0.045717f
C8346 AVDD.t17 AVSS 0.045717f
C8347 AVDD.n824 AVSS 0.537731f
C8348 AVDD.n825 AVSS 0.378581f
C8349 AVDD.n826 AVSS 0.712338f
C8350 AVDD.t450 AVSS 0.045717f
C8351 AVDD.t42 AVSS 0.045717f
C8352 AVDD.n827 AVSS 0.587661f
C8353 AVDD.t41 AVSS 0.089409f
C8354 AVDD.t449 AVSS 0.089409f
C8355 AVDD.n828 AVSS 0.445699f
C8356 AVDD.t700 AVSS 0.089409f
C8357 AVDD.t1017 AVSS 0.089409f
C8358 AVDD.n829 AVSS 0.445699f
C8359 AVDD.t1018 AVSS 0.045717f
C8360 AVDD.t701 AVSS 0.045717f
C8361 AVDD.n830 AVSS 0.764636f
C8362 AVDD.t573 AVSS 0.089409f
C8363 AVDD.t447 AVSS 0.089409f
C8364 AVDD.n831 AVSS 0.787444f
C8365 AVDD.t448 AVSS 0.045717f
C8366 AVDD.t574 AVSS 0.045717f
C8367 AVDD.n832 AVSS 0.446747f
C8368 AVDD.n833 AVSS 0.763137f
C8369 AVDD.t878 AVSS 0.045717f
C8370 AVDD.t978 AVSS 0.045717f
C8371 AVDD.n834 AVSS 0.446192f
C8372 AVDD.t977 AVSS 0.089409f
C8373 AVDD.t877 AVSS 0.089409f
C8374 AVDD.n835 AVSS 0.787444f
C8375 AVDD.t303 AVSS 0.045717f
C8376 AVDD.t397 AVSS 0.045717f
C8377 AVDD.n836 AVSS 0.764636f
C8378 AVDD.t396 AVSS 0.089409f
C8379 AVDD.t302 AVSS 0.089409f
C8380 AVDD.n837 AVSS 0.445699f
C8381 AVDD.t512 AVSS 0.089409f
C8382 AVDD.t401 AVSS 0.089409f
C8383 AVDD.n838 AVSS 0.445699f
C8384 AVDD.t402 AVSS 0.045717f
C8385 AVDD.t513 AVSS 0.045717f
C8386 AVDD.n839 AVSS 0.537731f
C8387 AVDD.n840 AVSS 0.712338f
C8388 AVDD.t386 AVSS 0.045717f
C8389 AVDD.t493 AVSS 0.045717f
C8390 AVDD.n841 AVSS 0.587661f
C8391 AVDD.t492 AVSS 0.089409f
C8392 AVDD.t385 AVSS 0.089409f
C8393 AVDD.n842 AVSS 0.445699f
C8394 AVDD.t613 AVSS 0.089409f
C8395 AVDD.t496 AVSS 0.089409f
C8396 AVDD.n843 AVSS 0.445699f
C8397 AVDD.t497 AVSS 0.045717f
C8398 AVDD.t614 AVSS 0.045717f
C8399 AVDD.n844 AVSS 0.743554f
C8400 AVDD.n845 AVSS 0.868895f
C8401 AVDD.t476 AVSS 0.033572f
C8402 AVDD.t76 AVSS 0.089409f
C8403 AVDD.n846 AVSS 0.363872f
C8404 AVDD.t961 AVSS 0.089409f
C8405 AVDD.n847 AVSS 0.340501f
C8406 AVDD.n848 AVSS 0.342168f
C8407 AVDD.t1260 AVSS 0.021426f
C8408 AVDD.t1005 AVSS 0.089409f
C8409 AVDD.n849 AVSS 0.173626f
C8410 AVDD.t1041 AVSS 0.089409f
C8411 AVDD.n850 AVSS 0.173626f
C8412 AVDD.n851 AVSS 0.141621f
C8413 AVDD.n852 AVSS 0.021426f
C8414 AVDD.t1042 AVSS 0.033572f
C8415 AVDD.n853 AVSS 0.148431f
C8416 AVDD.n854 AVSS 0.148431f
C8417 AVDD.t1006 AVSS 0.033572f
C8418 AVDD.n855 AVSS 0.021426f
C8419 AVDD.n856 AVSS 0.141621f
C8420 AVDD.t1259 AVSS 0.089409f
C8421 AVDD.n857 AVSS 0.173626f
C8422 AVDD.t616 AVSS 0.045717f
C8423 AVDD.n858 AVSS 0.245178f
C8424 AVDD.t879 AVSS 0.089409f
C8425 AVDD.n859 AVSS 0.473902f
C8426 AVDD.n860 AVSS 0.211727f
C8427 AVDD.n861 AVSS 0.021426f
C8428 AVDD.t880 AVSS 0.021426f
C8429 AVDD.t1153 AVSS 0.089409f
C8430 AVDD.n862 AVSS 0.363872f
C8431 AVDD.t615 AVSS 0.089409f
C8432 AVDD.n863 AVSS 0.363872f
C8433 AVDD.n864 AVSS 0.122697f
C8434 AVDD.n865 AVSS 0.021426f
C8435 AVDD.t1154 AVSS 0.033572f
C8436 AVDD.n866 AVSS 0.392415f
C8437 AVDD.n867 AVSS 0.392415f
C8438 AVDD.t475 AVSS 0.089409f
C8439 AVDD.n868 AVSS 0.363872f
C8440 AVDD.n869 AVSS 0.342168f
C8441 AVDD.t77 AVSS 0.045717f
C8442 AVDD.n870 AVSS 0.342168f
C8443 AVDD.n871 AVSS 0.331867f
C8444 AVDD.n872 AVSS 0.021426f
C8445 AVDD.t962 AVSS 0.021426f
C8446 AVDD.n873 AVSS 0.021426f
C8447 AVDD.n874 AVSS 0.308496f
C8448 AVDD.t901 AVSS 0.089409f
C8449 AVDD.n875 AVSS 0.363872f
C8450 AVDD.n876 AVSS 0.342168f
C8451 AVDD.t1250 AVSS 0.045717f
C8452 AVDD.n877 AVSS 0.342168f
C8453 AVDD.n878 AVSS 0.331867f
C8454 AVDD.n879 AVSS 0.021426f
C8455 AVDD.t687 AVSS 0.033572f
C8456 AVDD.n880 AVSS 0.342167f
C8457 AVDD.n881 AVSS 0.342167f
C8458 AVDD.t229 AVSS 0.033572f
C8459 AVDD.n882 AVSS 0.021426f
C8460 AVDD.n883 AVSS 0.331867f
C8461 AVDD.n884 AVSS 0.342167f
C8462 AVDD.t28 AVSS 0.033572f
C8463 AVDD.n885 AVSS 0.021426f
C8464 AVDD.t1122 AVSS 0.021426f
C8465 AVDD.n886 AVSS 0.021426f
C8466 AVDD.t1044 AVSS 0.033572f
C8467 AVDD.n887 AVSS 0.331651f
C8468 AVDD.t510 AVSS 0.089409f
C8469 AVDD.n888 AVSS 0.363872f
C8470 AVDD.t1043 AVSS 0.089409f
C8471 AVDD.n889 AVSS 0.363872f
C8472 AVDD.n890 AVSS 0.331867f
C8473 AVDD.n891 AVSS 0.021426f
C8474 AVDD.t65 AVSS 0.021426f
C8475 AVDD.n892 AVSS 0.021426f
C8476 AVDD.n893 AVSS 0.045573f
C8477 AVDD.n894 AVSS 0.326024f
C8478 AVDD.n895 AVSS 0.416263f
C8479 AVDD.n896 AVSS 0.417334f
C8480 AVDD.t13 AVSS 4.59466f
C8481 AVDD.n897 AVSS 0.206501f
C8482 AVDD.n898 AVSS 0.207284f
C8483 AVDD.t783 AVSS 0.089409f
C8484 AVDD.n899 AVSS 0.190118f
C8485 AVDD.t784 AVSS 0.045717f
C8486 AVDD.t1150 AVSS 0.026723f
C8487 AVDD.t805 AVSS 0.058154f
C8488 AVDD.n900 AVSS 0.239368f
C8489 AVDD.n901 AVSS 0.006326f
C8490 AVDD.t1695 AVSS 0.010713f
C8491 AVDD.t1601 AVSS 0.010713f
C8492 AVDD.n902 AVSS 0.024453f
C8493 AVDD.n903 AVSS 0.021084f
C8494 AVDD.n904 AVSS 0.006326f
C8495 AVDD.t1598 AVSS 0.010713f
C8496 AVDD.t1698 AVSS 0.010713f
C8497 AVDD.n905 AVSS 0.024453f
C8498 AVDD.n906 AVSS 0.021084f
C8499 AVDD.n907 AVSS 0.006326f
C8500 AVDD.t1427 AVSS 0.025859f
C8501 AVDD.n908 AVSS 0.031411f
C8502 AVDD.n909 AVSS 0.006326f
C8503 AVDD.t1650 AVSS 0.010713f
C8504 AVDD.t1587 AVSS 0.010713f
C8505 AVDD.n910 AVSS 0.024453f
C8506 AVDD.n911 AVSS 0.021084f
C8507 AVDD.n912 AVSS 0.006326f
C8508 AVDD.t1283 AVSS 0.010713f
C8509 AVDD.t1693 AVSS 0.010713f
C8510 AVDD.n913 AVSS 0.024453f
C8511 AVDD.n914 AVSS 0.021084f
C8512 AVDD.n915 AVSS 0.006326f
C8513 AVDD.t1699 AVSS 0.010713f
C8514 AVDD.t1281 AVSS 0.010713f
C8515 AVDD.n916 AVSS 0.024453f
C8516 AVDD.n917 AVSS 0.021084f
C8517 AVDD.t817 AVSS 0.045717f
C8518 AVDD.n918 AVSS 0.198115f
C8519 AVDD.t246 AVSS 0.045717f
C8520 AVDD.t809 AVSS 0.089409f
C8521 AVDD.n919 AVSS 0.169461f
C8522 AVDD.t324 AVSS 0.021426f
C8523 AVDD.t1221 AVSS 0.089409f
C8524 AVDD.n920 AVSS 0.169461f
C8525 AVDD.t876 AVSS 0.033572f
C8526 AVDD.t637 AVSS 0.089409f
C8527 AVDD.n921 AVSS 0.169461f
C8528 AVDD.t718 AVSS 0.021426f
C8529 AVDD.t925 AVSS 0.089409f
C8530 AVDD.n922 AVSS 0.169461f
C8531 AVDD.t281 AVSS 0.089409f
C8532 AVDD.n923 AVSS 0.169461f
C8533 AVDD.t481 AVSS 0.021426f
C8534 AVDD.t554 AVSS 0.089409f
C8535 AVDD.n924 AVSS 0.169461f
C8536 AVDD.t40 AVSS 0.033572f
C8537 AVDD.t806 AVSS 0.026723f
C8538 AVDD.n925 AVSS 0.277143f
C8539 AVDD.t190 AVSS 0.089409f
C8540 AVDD.n926 AVSS 0.263904f
C8541 AVDD.t387 AVSS 0.058154f
C8542 AVDD.n927 AVSS 0.187773f
C8543 AVDD.t191 AVSS 0.045717f
C8544 AVDD.n928 AVSS 0.121571f
C8545 AVDD.t388 AVSS 0.026723f
C8546 AVDD.t666 AVSS 0.058154f
C8547 AVDD.n929 AVSS 0.12966f
C8548 AVDD.t742 AVSS 0.012856f
C8549 AVDD.n930 AVSS 0.053606f
C8550 AVDD.t1379 AVSS 0.015123f
C8551 AVDD.t991 AVSS 0.058154f
C8552 AVDD.n931 AVSS 0.130566f
C8553 AVDD.t1183 AVSS 0.058154f
C8554 AVDD.n932 AVSS 0.108676f
C8555 AVDD.t395 AVSS 0.012856f
C8556 AVDD.n933 AVSS 0.054058f
C8557 AVDD.t327 AVSS 0.058154f
C8558 AVDD.n934 AVSS 0.130566f
C8559 AVDD.t14 AVSS 0.026723f
C8560 AVDD.t932 AVSS 0.026723f
C8561 AVDD.t659 AVSS 0.045717f
C8562 AVDD.t898 AVSS 0.026723f
C8563 AVDD.n935 AVSS 0.229432f
C8564 AVDD.t658 AVSS 0.089409f
C8565 AVDD.n936 AVSS 0.152947f
C8566 AVDD.t897 AVSS 0.058154f
C8567 AVDD.n937 AVSS 0.187773f
C8568 AVDD.n938 AVSS 0.180933f
C8569 AVDD.t931 AVSS 0.058154f
C8570 AVDD.n939 AVSS 0.189993f
C8571 AVDD.n940 AVSS 0.166742f
C8572 AVDD.t1142 AVSS 0.045717f
C8573 AVDD.n941 AVSS 0.230095f
C8574 AVDD.t1141 AVSS 0.089409f
C8575 AVDD.n942 AVSS 0.20708f
C8576 AVDD.t707 AVSS 0.045717f
C8577 AVDD.t816 AVSS 0.089409f
C8578 AVDD.n943 AVSS 0.218463f
C8579 AVDD.t706 AVSS 0.089409f
C8580 AVDD.n944 AVSS 0.218463f
C8581 AVDD.n945 AVSS 0.199199f
C8582 AVDD.n946 AVSS 0.208268f
C8583 AVDD.t1291 AVSS 0.010713f
C8584 AVDD.t1653 AVSS 0.010713f
C8585 AVDD.n947 AVSS 0.038647f
C8586 AVDD.n948 AVSS 0.096508f
C8587 AVDD.t1640 AVSS 0.010713f
C8588 AVDD.t1384 AVSS 0.010713f
C8589 AVDD.n949 AVSS 0.038647f
C8590 AVDD.n950 AVSS 0.071452f
C8591 AVDD.t1685 AVSS 0.038924f
C8592 AVDD.n951 AVSS 0.082909f
C8593 AVDD.t1415 AVSS 0.010713f
C8594 AVDD.t1676 AVSS 0.010713f
C8595 AVDD.n952 AVSS 0.038647f
C8596 AVDD.n953 AVSS 0.085941f
C8597 AVDD.t1576 AVSS 0.010713f
C8598 AVDD.t1461 AVSS 0.010713f
C8599 AVDD.n954 AVSS 0.038647f
C8600 AVDD.n955 AVSS 0.08594f
C8601 AVDD.t1457 AVSS 0.010713f
C8602 AVDD.t1568 AVSS 0.010713f
C8603 AVDD.n956 AVSS 0.038647f
C8604 AVDD.n957 AVSS 0.096235f
C8605 AVDD.n958 AVSS 0.241665f
C8606 AVDD.t1079 AVSS 0.089409f
C8607 AVDD.n959 AVSS 0.231171f
C8608 AVDD.t12 AVSS 0.058154f
C8609 AVDD.n960 AVSS 0.149494f
C8610 AVDD.n961 AVSS 0.157311f
C8611 AVDD.n962 AVSS 0.09329f
C8612 AVDD.n963 AVSS 0.115602f
C8613 AVDD.t329 AVSS 0.019789f
C8614 AVDD.n964 AVSS 0.012856f
C8615 AVDD.n965 AVSS 0.108117f
C8616 AVDD.t393 AVSS 0.058154f
C8617 AVDD.n966 AVSS 0.130566f
C8618 AVDD.n967 AVSS 0.075948f
C8619 AVDD.n968 AVSS 0.012856f
C8620 AVDD.t1184 AVSS 0.019789f
C8621 AVDD.n969 AVSS 0.111605f
C8622 AVDD.n970 AVSS 0.111605f
C8623 AVDD.t992 AVSS 0.026723f
C8624 AVDD.n971 AVSS 0.131878f
C8625 AVDD.t1276 AVSS 0.026723f
C8626 AVDD.n972 AVSS 0.283157f
C8627 AVDD.t1275 AVSS 0.058154f
C8628 AVDD.n973 AVSS 0.195624f
C8629 AVDD.t920 AVSS 0.026723f
C8630 AVDD.n974 AVSS 0.186243f
C8631 AVDD.t919 AVSS 0.058154f
C8632 AVDD.n975 AVSS 0.156405f
C8633 AVDD.t887 AVSS 0.058154f
C8634 AVDD.t542 AVSS 0.058154f
C8635 AVDD.n976 AVSS 0.267564f
C8636 AVDD.t543 AVSS 0.026723f
C8637 AVDD.t888 AVSS 0.026723f
C8638 AVDD.n977 AVSS 0.30086f
C8639 AVDD.t328 AVSS 4.90298f
C8640 AVDD.t394 AVSS 3.24073f
C8641 AVDD.n978 AVSS 1.90355f
C8642 AVDD.t264 AVSS 3.36808f
C8643 AVDD.t2 AVSS 5.68049f
C8644 AVDD.t373 AVSS 4.48225f
C8645 AVDD.n979 AVSS 2.45788f
C8646 AVDD.n980 AVSS 0.320056f
C8647 AVDD.t808 AVSS 0.026723f
C8648 AVDD.t1132 AVSS 0.026723f
C8649 AVDD.n981 AVSS 0.309598f
C8650 AVDD.t1131 AVSS 0.058154f
C8651 AVDD.t807 AVSS 0.058154f
C8652 AVDD.n982 AVSS 0.321806f
C8653 AVDD.t797 AVSS 0.058154f
C8654 AVDD.t435 AVSS 0.058154f
C8655 AVDD.n983 AVSS 0.321806f
C8656 AVDD.t436 AVSS 0.026723f
C8657 AVDD.t798 AVSS 0.026723f
C8658 AVDD.n984 AVSS 0.373501f
C8659 AVDD.t372 AVSS 0.058154f
C8660 AVDD.t1 AVSS 0.058154f
C8661 AVDD.n985 AVSS 0.275928f
C8662 AVDD.t3 AVSS 0.026723f
C8663 AVDD.t374 AVSS 0.026723f
C8664 AVDD.n986 AVSS 0.509497f
C8665 AVDD.n987 AVSS 0.236032f
C8666 AVDD.t263 AVSS 0.058154f
C8667 AVDD.n988 AVSS 0.127323f
C8668 AVDD.n989 AVSS 0.102048f
C8669 AVDD.t265 AVSS 0.019789f
C8670 AVDD.n990 AVSS 0.012856f
C8671 AVDD.n991 AVSS 0.075312f
C8672 AVDD.t741 AVSS 0.058154f
C8673 AVDD.n992 AVSS 0.12966f
C8674 AVDD.n993 AVSS 0.107212f
C8675 AVDD.n994 AVSS 0.012856f
C8676 AVDD.t667 AVSS 0.019789f
C8677 AVDD.n995 AVSS 0.13326f
C8678 AVDD.n996 AVSS 0.449598f
C8679 AVDD.n997 AVSS 0.11432f
C8680 AVDD.n998 AVSS 0.148966f
C8681 AVDD.t38 AVSS 0.089409f
C8682 AVDD.n999 AVSS 0.169461f
C8683 AVDD.n1000 AVSS 0.137456f
C8684 AVDD.n1001 AVSS 0.021426f
C8685 AVDD.t556 AVSS 0.021426f
C8686 AVDD.n1002 AVSS 0.021426f
C8687 AVDD.n1003 AVSS 0.137456f
C8688 AVDD.t479 AVSS 0.089409f
C8689 AVDD.n1004 AVSS 0.169461f
C8690 AVDD.n1005 AVSS 0.137456f
C8691 AVDD.n1006 AVSS 0.021426f
C8692 AVDD.t283 AVSS 0.033572f
C8693 AVDD.n1007 AVSS 0.144368f
C8694 AVDD.n1008 AVSS 0.144368f
C8695 AVDD.t926 AVSS 0.033572f
C8696 AVDD.n1009 AVSS 0.021426f
C8697 AVDD.n1010 AVSS 0.128017f
C8698 AVDD.n1011 AVSS 0.068727f
C8699 AVDD.t716 AVSS 0.089409f
C8700 AVDD.n1012 AVSS 0.110171f
C8701 AVDD.n1013 AVSS 0.137456f
C8702 AVDD.n1014 AVSS 0.021426f
C8703 AVDD.t639 AVSS 0.033572f
C8704 AVDD.n1015 AVSS 0.144368f
C8705 AVDD.n1016 AVSS 0.144368f
C8706 AVDD.t874 AVSS 0.089409f
C8707 AVDD.n1017 AVSS 0.169461f
C8708 AVDD.n1018 AVSS 0.137456f
C8709 AVDD.n1019 AVSS 0.021426f
C8710 AVDD.t1222 AVSS 0.021426f
C8711 AVDD.n1020 AVSS 0.021426f
C8712 AVDD.n1021 AVSS 0.137456f
C8713 AVDD.t322 AVSS 0.089409f
C8714 AVDD.n1022 AVSS 0.169461f
C8715 AVDD.n1023 AVSS 0.137456f
C8716 AVDD.n1024 AVSS 0.021426f
C8717 AVDD.t811 AVSS 0.033572f
C8718 AVDD.n1025 AVSS 0.183348f
C8719 AVDD.n1026 AVSS 0.366195f
C8720 AVDD.t245 AVSS 0.089409f
C8721 AVDD.n1027 AVSS 0.288655f
C8722 AVDD.n1028 AVSS 0.286344f
C8723 AVDD.n1029 AVSS 0.046036f
C8724 AVDD.n1030 AVSS 0.014056f
C8725 AVDD.n1031 AVSS 0.025912f
C8726 AVDD.n1032 AVSS 0.025919f
C8727 AVDD.n1033 AVSS 0.014056f
C8728 AVDD.n1034 AVSS 0.032799f
C8729 AVDD.n1035 AVSS 0.032805f
C8730 AVDD.n1036 AVSS 0.014056f
C8731 AVDD.n1037 AVSS 0.025912f
C8732 AVDD.n1038 AVSS 0.025919f
C8733 AVDD.n1039 AVSS 0.014056f
C8734 AVDD.n1040 AVSS 0.018311f
C8735 AVDD.n1041 AVSS 0.018317f
C8736 AVDD.n1042 AVSS 0.014056f
C8737 AVDD.n1043 AVSS 0.025912f
C8738 AVDD.n1044 AVSS 0.025919f
C8739 AVDD.n1045 AVSS 0.014056f
C8740 AVDD.n1046 AVSS 0.045772f
C8741 AVDD.n1047 AVSS 0.173835f
C8742 AVDD.t1149 AVSS 0.058154f
C8743 AVDD.n1048 AVSS 0.207745f
C8744 AVDD.n1049 AVSS 0.14677f
C8745 AVDD.n1050 AVSS 0.18759f
C8746 AVDD.n1051 AVSS 0.165325f
C8747 AVDD.n1052 AVSS 0.207229f
C8748 AVDD.n1053 AVSS 2.07782f
C8749 AVDD.n1054 AVSS 17.6971f
C8750 AVDD.t181 AVSS 4.62261f
C8751 AVDD.t810 AVSS 4.90298f
C8752 AVDD.t323 AVSS 3.8071f
C8753 AVDD.t366 AVSS 3.8071f
C8754 AVDD.t875 AVSS 4.71196f
C8755 AVDD.t638 AVSS 4.71196f
C8756 AVDD.t717 AVSS 2.03425f
C8757 AVDD.n1055 AVSS 1.90355f
C8758 AVDD.t27 AVSS 4.1858f
C8759 AVDD.t33 AVSS 13.1202f
C8760 AVDD.t85 AVSS 10.1876f
C8761 AVDD.t378 AVSS 10.1876f
C8762 AVDD.t93 AVSS 12.609f
C8763 AVDD.t233 AVSS 12.609f
C8764 AVDD.t186 AVSS 5.3808f
C8765 AVDD.n1056 AVSS 5.09382f
C8766 AVDD.t238 AVSS 12.322001f
C8767 AVDD.t82 AVSS 12.609f
C8768 AVDD.t36 AVSS 10.1876f
C8769 AVDD.t255 AVSS 10.1876f
C8770 AVDD.t205 AVSS 8.95903f
C8771 AVDD.n1057 AVSS 10.8348f
C8772 AVDD.t282 AVSS 2.29901f
C8773 AVDD.t480 AVSS 3.8071f
C8774 AVDD.t555 AVSS 3.8071f
C8775 AVDD.t39 AVSS 4.90298f
C8776 AVDD.t131 AVSS 4.59466f
C8777 AVDD.n1058 AVSS 2.07782f
C8778 AVDD.n1059 AVSS 0.415071f
C8779 AVDD.n1060 AVSS 0.15613f
C8780 AVDD.n1061 AVSS 0.14196f
C8781 AVDD.n1062 AVSS 0.045683f
C8782 AVDD.t1455 AVSS 0.010713f
C8783 AVDD.t1565 AVSS 0.010713f
C8784 AVDD.n1063 AVSS 0.025023f
C8785 AVDD.n1064 AVSS 0.02284f
C8786 AVDD.t1574 AVSS 0.010713f
C8787 AVDD.t1436 AVSS 0.010713f
C8788 AVDD.n1065 AVSS 0.026795f
C8789 AVDD.n1066 AVSS 0.039995f
C8790 AVDD.n1067 AVSS 0.025919f
C8791 AVDD.n1068 AVSS 0.025912f
C8792 AVDD.t1575 AVSS 0.010713f
C8793 AVDD.t1302 AVSS 0.010713f
C8794 AVDD.n1069 AVSS 0.025023f
C8795 AVDD.n1070 AVSS 0.02284f
C8796 AVDD.t1418 AVSS 0.010713f
C8797 AVDD.t1677 AVSS 0.010713f
C8798 AVDD.n1071 AVSS 0.026795f
C8799 AVDD.n1072 AVSS 0.039995f
C8800 AVDD.n1073 AVSS 0.018317f
C8801 AVDD.n1074 AVSS 0.018311f
C8802 AVDD.t1282 AVSS 0.026362f
C8803 AVDD.n1075 AVSS 0.033235f
C8804 AVDD.t1694 AVSS 0.027891f
C8805 AVDD.n1076 AVSS 0.050632f
C8806 AVDD.n1077 AVSS 0.025919f
C8807 AVDD.n1078 AVSS 0.025912f
C8808 AVDD.t1602 AVSS 0.010713f
C8809 AVDD.t1600 AVSS 0.010713f
C8810 AVDD.n1079 AVSS 0.025023f
C8811 AVDD.n1080 AVSS 0.02284f
C8812 AVDD.t1692 AVSS 0.010713f
C8813 AVDD.t1284 AVSS 0.010713f
C8814 AVDD.n1081 AVSS 0.026795f
C8815 AVDD.n1082 AVSS 0.039995f
C8816 AVDD.n1083 AVSS 0.032805f
C8817 AVDD.n1084 AVSS 0.032799f
C8818 AVDD.t1426 AVSS 0.010713f
C8819 AVDD.t1381 AVSS 0.010713f
C8820 AVDD.n1085 AVSS 0.025023f
C8821 AVDD.n1086 AVSS 0.02284f
C8822 AVDD.t1486 AVSS 0.010713f
C8823 AVDD.t1666 AVSS 0.010713f
C8824 AVDD.n1087 AVSS 0.026795f
C8825 AVDD.n1088 AVSS 0.039995f
C8826 AVDD.n1089 AVSS 0.025919f
C8827 AVDD.n1090 AVSS 0.025912f
C8828 AVDD.t1290 AVSS 0.010713f
C8829 AVDD.t1651 AVSS 0.010713f
C8830 AVDD.n1091 AVSS 0.025023f
C8831 AVDD.n1092 AVSS 0.02284f
C8832 AVDD.t1585 AVSS 0.010713f
C8833 AVDD.t1382 AVSS 0.010713f
C8834 AVDD.n1093 AVSS 0.026795f
C8835 AVDD.n1094 AVSS 0.039995f
C8836 AVDD.n1095 AVSS 0.046066f
C8837 AVDD.n1096 AVSS 0.141644f
C8838 AVDD.n1097 AVSS 0.210311f
C8839 AVDD.t723 AVSS 0.089409f
C8840 AVDD.n1098 AVSS 0.206538f
C8841 AVDD.n1099 AVSS 0.200663f
C8842 AVDD.n1100 AVSS 0.045977f
C8843 AVDD.n1101 AVSS 0.014057f
C8844 AVDD.n1102 AVSS 0.025911f
C8845 AVDD.n1103 AVSS 0.02592f
C8846 AVDD.n1104 AVSS 0.014057f
C8847 AVDD.n1105 AVSS 0.032798f
C8848 AVDD.n1106 AVSS 0.032807f
C8849 AVDD.n1107 AVSS 0.014057f
C8850 AVDD.n1108 AVSS 0.025911f
C8851 AVDD.n1109 AVSS 0.02592f
C8852 AVDD.n1110 AVSS 0.014057f
C8853 AVDD.n1111 AVSS 0.01831f
C8854 AVDD.n1112 AVSS 0.018319f
C8855 AVDD.n1113 AVSS 0.014057f
C8856 AVDD.n1114 AVSS 0.025911f
C8857 AVDD.n1115 AVSS 0.02592f
C8858 AVDD.n1116 AVSS 0.014057f
C8859 AVDD.n1117 AVSS 0.045713f
C8860 AVDD.n1118 AVSS 0.201338f
C8861 AVDD.n1119 AVSS 0.195411f
C8862 AVDD.t130 AVSS 0.089409f
C8863 AVDD.n1120 AVSS 0.21934f
C8864 AVDD.t945 AVSS 0.089409f
C8865 AVDD.n1121 AVSS 0.21934f
C8866 AVDD.n1122 AVSS 0.207391f
C8867 AVDD.n1123 AVSS 0.279517f
C8868 AVDD.t1697 AVSS 0.010713f
C8869 AVDD.t1604 AVSS 0.010713f
C8870 AVDD.n1124 AVSS 0.039216f
C8871 AVDD.n1125 AVSS 0.097035f
C8872 AVDD.t1603 AVSS 0.010713f
C8873 AVDD.t1597 AVSS 0.010713f
C8874 AVDD.n1126 AVSS 0.039216f
C8875 AVDD.n1127 AVSS 0.086657f
C8876 AVDD.t1390 AVSS 0.010713f
C8877 AVDD.t1434 AVSS 0.010713f
C8878 AVDD.n1128 AVSS 0.039303f
C8879 AVDD.n1129 AVSS 0.086739f
C8880 AVDD.t1414 AVSS 0.039472f
C8881 AVDD.n1130 AVSS 0.083816f
C8882 AVDD.t1691 AVSS 0.010713f
C8883 AVDD.t1696 AVSS 0.010713f
C8884 AVDD.n1131 AVSS 0.039216f
C8885 AVDD.n1132 AVSS 0.072168f
C8886 AVDD.t1599 AVSS 0.010713f
C8887 AVDD.t1285 AVSS 0.010713f
C8888 AVDD.n1133 AVSS 0.039216f
C8889 AVDD.n1134 AVSS 0.097365f
C8890 AVDD.n1135 AVSS 0.278577f
C8891 AVDD.t1185 AVSS 0.089409f
C8892 AVDD.n1136 AVSS 0.243512f
C8893 AVDD.n1137 AVSS 0.416605f
C8894 AVDD.t654 AVSS 0.089409f
C8895 AVDD.n1138 AVSS 0.224815f
C8896 AVDD.n1139 AVSS 0.331867f
C8897 AVDD.n1140 AVSS 0.021426f
C8898 AVDD.t1186 AVSS 0.021426f
C8899 AVDD.n1141 AVSS 0.021426f
C8900 AVDD.n1142 AVSS 0.374556f
C8901 AVDD.t789 AVSS 0.089409f
C8902 AVDD.n1143 AVSS 0.169743f
C8903 AVDD.n1144 AVSS 0.141621f
C8904 AVDD.n1145 AVSS 0.021426f
C8905 AVDD.t740 AVSS 0.033572f
C8906 AVDD.n1146 AVSS 0.197655f
C8907 AVDD.n1147 AVSS 0.374471f
C8908 AVDD.t1261 AVSS 0.089409f
C8909 AVDD.n1148 AVSS 0.389564f
C8910 AVDD.n1149 AVSS 0.37816f
C8911 AVDD.t516 AVSS 0.089409f
C8912 AVDD.n1150 AVSS 0.220656f
C8913 AVDD.t405 AVSS 0.089409f
C8914 AVDD.n1151 AVSS 0.220656f
C8915 AVDD.n1152 AVSS 0.29069f
C8916 AVDD.n1153 AVSS 0.352075f
C8917 AVDD.n1154 AVSS 0.378581f
C8918 AVDD.t61 AVSS 0.089409f
C8919 AVDD.n1155 AVSS 0.389564f
C8920 AVDD.t596 AVSS 0.045717f
C8921 AVDD.n1156 AVSS 0.37816f
C8922 AVDD.t595 AVSS 0.089409f
C8923 AVDD.n1157 AVSS 0.220656f
C8924 AVDD.t486 AVSS 0.089409f
C8925 AVDD.n1158 AVSS 0.220656f
C8926 AVDD.t487 AVSS 0.045717f
C8927 AVDD.n1159 AVSS 0.266012f
C8928 AVDD.t564 AVSS 0.045717f
C8929 AVDD.t776 AVSS 0.045717f
C8930 AVDD.t621 AVSS 0.089409f
C8931 AVDD.t1245 AVSS 0.089409f
C8932 AVDD.n1160 AVSS 0.256112f
C8933 AVDD.t622 AVSS 0.045717f
C8934 AVDD.t32 AVSS 0.089409f
C8935 AVDD.t714 AVSS 0.089409f
C8936 AVDD.n1161 AVSS 0.342362f
C8937 AVDD.t34 AVSS 0.033572f
C8938 AVDD.t766 AVSS 0.021426f
C8939 AVDD.t84 AVSS 0.089409f
C8940 AVDD.t765 AVSS 0.089409f
C8941 AVDD.n1162 AVSS 0.342362f
C8942 AVDD.t519 AVSS 0.021426f
C8943 AVDD.t518 AVSS 0.089409f
C8944 AVDD.t1169 AVSS 0.089409f
C8945 AVDD.n1163 AVSS 0.342362f
C8946 AVDD.t900 AVSS 0.033572f
C8947 AVDD.t257 AVSS 0.089409f
C8948 AVDD.t899 AVSS 0.089409f
C8949 AVDD.n1164 AVSS 0.342362f
C8950 AVDD.t1239 AVSS 0.089409f
C8951 AVDD.t619 AVSS 0.089409f
C8952 AVDD.n1165 AVSS 0.342362f
C8953 AVDD.t1240 AVSS 0.033572f
C8954 AVDD.t187 AVSS 0.021426f
C8955 AVDD.t840 AVSS 0.089409f
C8956 AVDD.t185 AVSS 0.089409f
C8957 AVDD.n1166 AVSS 0.218868f
C8958 AVDD.t884 AVSS 0.033572f
C8959 AVDD.t883 AVSS 0.089409f
C8960 AVDD.t237 AVSS 0.089409f
C8961 AVDD.n1167 AVSS 0.342362f
C8962 AVDD.n1168 AVSS 0.139176f
C8963 AVDD.t1113 AVSS 0.089409f
C8964 AVDD.t488 AVSS 0.089409f
C8965 AVDD.n1169 AVSS 0.342362f
C8966 AVDD.t1114 AVSS 0.033572f
C8967 AVDD.t37 AVSS 0.021426f
C8968 AVDD.t704 AVSS 0.089409f
C8969 AVDD.t35 AVSS 0.089409f
C8970 AVDD.n1170 AVSS 0.342362f
C8971 AVDD.t1244 AVSS 0.021426f
C8972 AVDD.t1243 AVSS 0.089409f
C8973 AVDD.t627 AVSS 0.089409f
C8974 AVDD.n1171 AVSS 0.342362f
C8975 AVDD.t206 AVSS 0.033572f
C8976 AVDD.t850 AVSS 0.089409f
C8977 AVDD.t204 AVSS 0.089409f
C8978 AVDD.n1172 AVSS 0.342362f
C8979 AVDD.t851 AVSS 0.033572f
C8980 AVDD.n1173 AVSS 0.021426f
C8981 AVDD.n1174 AVSS 0.278352f
C8982 AVDD.n1175 AVSS 0.021426f
C8983 AVDD.t628 AVSS 0.021426f
C8984 AVDD.n1176 AVSS 0.021426f
C8985 AVDD.n1177 AVSS 0.278352f
C8986 AVDD.n1178 AVSS 0.021426f
C8987 AVDD.t705 AVSS 0.021426f
C8988 AVDD.n1179 AVSS 0.021426f
C8989 AVDD.n1180 AVSS 0.278352f
C8990 AVDD.n1181 AVSS 0.021426f
C8991 AVDD.t489 AVSS 0.033572f
C8992 AVDD.n1182 AVSS 0.292092f
C8993 AVDD.n1183 AVSS 0.292092f
C8994 AVDD.t239 AVSS 0.033572f
C8995 AVDD.n1184 AVSS 0.021426f
C8996 AVDD.n1185 AVSS 0.26267f
C8997 AVDD.n1186 AVSS 0.021426f
C8998 AVDD.t841 AVSS 0.021426f
C8999 AVDD.n1187 AVSS 0.021426f
C9000 AVDD.n1188 AVSS 0.278352f
C9001 AVDD.n1189 AVSS 0.021426f
C9002 AVDD.t620 AVSS 0.033572f
C9003 AVDD.n1190 AVSS 0.292092f
C9004 AVDD.n1191 AVSS 0.292092f
C9005 AVDD.t258 AVSS 0.033572f
C9006 AVDD.n1192 AVSS 0.021426f
C9007 AVDD.n1193 AVSS 0.278352f
C9008 AVDD.n1194 AVSS 0.021426f
C9009 AVDD.t1170 AVSS 0.021426f
C9010 AVDD.n1195 AVSS 0.021426f
C9011 AVDD.n1196 AVSS 0.278352f
C9012 AVDD.n1197 AVSS 0.021426f
C9013 AVDD.t86 AVSS 0.021426f
C9014 AVDD.n1198 AVSS 0.021426f
C9015 AVDD.n1199 AVSS 0.278352f
C9016 AVDD.n1200 AVSS 0.021426f
C9017 AVDD.t715 AVSS 0.033572f
C9018 AVDD.n1201 AVSS 0.320025f
C9019 AVDD.n1202 AVSS 0.320025f
C9020 AVDD.t1246 AVSS 0.045717f
C9021 AVDD.n1203 AVSS 0.3558f
C9022 AVDD.t1130 AVSS 0.045717f
C9023 AVDD.t1014 AVSS 0.045717f
C9024 AVDD.t936 AVSS 0.045717f
C9025 AVDD.t832 AVSS 0.089409f
C9026 AVDD.n1204 AVSS 0.220656f
C9027 AVDD.t935 AVSS 0.089409f
C9028 AVDD.n1205 AVSS 0.220656f
C9029 AVDD.n1206 AVSS 0.29069f
C9030 AVDD.n1207 AVSS 0.352075f
C9031 AVDD.n1208 AVSS 0.266012f
C9032 AVDD.t1013 AVSS 0.089409f
C9033 AVDD.n1209 AVSS 0.220656f
C9034 AVDD.t1129 AVSS 0.089409f
C9035 AVDD.n1210 AVSS 0.220656f
C9036 AVDD.n1211 AVSS 0.367741f
C9037 AVDD.n1212 AVSS 0.670031f
C9038 AVDD.n1213 AVSS 0.367741f
C9039 AVDD.t775 AVSS 0.089409f
C9040 AVDD.n1214 AVSS 0.220656f
C9041 AVDD.t563 AVSS 0.089409f
C9042 AVDD.n1215 AVSS 0.220656f
C9043 AVDD.n1216 AVSS 0.29069f
C9044 AVDD.n1217 AVSS 0.352075f
C9045 AVDD.n1218 AVSS 0.378581f
C9046 AVDD.n1219 AVSS 5.90094f
C9047 AVDD.n1220 AVSS 0.378581f
C9048 AVDD.n1221 AVSS 0.352075f
C9049 AVDD.n1222 AVSS 0.266012f
C9050 AVDD.t514 AVSS 0.089409f
C9051 AVDD.n1223 AVSS 0.220656f
C9052 AVDD.t625 AVSS 0.089409f
C9053 AVDD.n1224 AVSS 0.220656f
C9054 AVDD.n1225 AVSS 0.367741f
C9055 AVDD.n1226 AVSS 0.775975f
C9056 AVDD.n1227 AVSS 0.61096f
C9057 AVDD.t105 AVSS 0.045717f
C9058 AVDD.n1228 AVSS 0.547954f
C9059 AVDD.n1229 AVSS 0.547954f
C9060 AVDD.t664 AVSS 0.089409f
C9061 AVDD.n1230 AVSS 0.55425f
C9062 AVDD.n1231 AVSS 0.49024f
C9063 AVDD.n1232 AVSS 0.021426f
C9064 AVDD.t285 AVSS 0.021426f
C9065 AVDD.n1233 AVSS 0.021426f
C9066 AVDD.n1234 AVSS 0.49024f
C9067 AVDD.t965 AVSS 0.089409f
C9068 AVDD.n1235 AVSS 0.55425f
C9069 AVDD.n1236 AVSS 0.49024f
C9070 AVDD.n1237 AVSS 0.021426f
C9071 AVDD.t904 AVSS 0.033572f
C9072 AVDD.n1238 AVSS 0.498758f
C9073 AVDD.n1239 AVSS 0.498758f
C9074 AVDD.t527 AVSS 0.033572f
C9075 AVDD.n1240 AVSS 0.021426f
C9076 AVDD.n1241 AVSS 0.49024f
C9077 AVDD.t905 AVSS 0.089409f
C9078 AVDD.n1242 AVSS 0.33675f
C9079 AVDD.n1243 AVSS 0.24512f
C9080 AVDD.n1244 AVSS 0.462621f
C9081 AVDD.n1245 AVSS 0.021426f
C9082 AVDD.t501 AVSS 0.033572f
C9083 AVDD.n1246 AVSS 0.498758f
C9084 AVDD.n1247 AVSS 0.498758f
C9085 AVDD.t90 AVSS 0.089409f
C9086 AVDD.n1248 AVSS 0.55425f
C9087 AVDD.n1249 AVSS 0.49024f
C9088 AVDD.n1250 AVSS 0.021426f
C9089 AVDD.t472 AVSS 0.021426f
C9090 AVDD.n1251 AVSS 0.021426f
C9091 AVDD.n1252 AVSS 0.49024f
C9092 AVDD.t747 AVSS 0.089409f
C9093 AVDD.n1253 AVSS 0.55425f
C9094 AVDD.n1254 AVSS 0.49024f
C9095 AVDD.n1255 AVSS 0.021426f
C9096 AVDD.t1098 AVSS 0.033572f
C9097 AVDD.n1256 AVSS 0.547954f
C9098 AVDD.n1257 AVSS 0.547954f
C9099 AVDD.t9 AVSS 0.045717f
C9100 AVDD.n1258 AVSS 0.493579f
C9101 AVDD.t457 AVSS 0.089409f
C9102 AVDD.t881 AVSS 0.089409f
C9103 AVDD.n1259 AVSS 0.445699f
C9104 AVDD.t357 AVSS 0.089409f
C9105 AVDD.t773 AVSS 0.089409f
C9106 AVDD.n1260 AVSS 0.445699f
C9107 AVDD.t774 AVSS 0.045717f
C9108 AVDD.t358 AVSS 0.045717f
C9109 AVDD.n1261 AVSS 0.743554f
C9110 AVDD.n1262 AVSS 1.52977f
C9111 AVDD.n1263 AVSS 0.493579f
C9112 AVDD.t938 AVSS 0.045717f
C9113 AVDD.n1264 AVSS 0.547954f
C9114 AVDD.n1265 AVSS 0.547954f
C9115 AVDD.t1157 AVSS 0.089409f
C9116 AVDD.n1266 AVSS 0.55425f
C9117 AVDD.n1267 AVSS 0.49024f
C9118 AVDD.n1268 AVSS 0.021426f
C9119 AVDD.t1068 AVSS 0.021426f
C9120 AVDD.n1269 AVSS 0.021426f
C9121 AVDD.n1270 AVSS 0.49024f
C9122 AVDD.t494 AVSS 0.089409f
C9123 AVDD.n1271 AVSS 0.55425f
C9124 AVDD.n1272 AVSS 0.49024f
C9125 AVDD.n1273 AVSS 0.021426f
C9126 AVDD.t426 AVSS 0.033572f
C9127 AVDD.n1274 AVSS 0.498758f
C9128 AVDD.n1275 AVSS 0.498758f
C9129 AVDD.t1016 AVSS 0.033572f
C9130 AVDD.n1276 AVSS 0.021426f
C9131 AVDD.n1277 AVSS 0.49024f
C9132 AVDD.t97 AVSS 0.089409f
C9133 AVDD.n1278 AVSS 0.33675f
C9134 AVDD.n1279 AVSS 0.24512f
C9135 AVDD.n1280 AVSS 0.462621f
C9136 AVDD.n1281 AVSS 0.021426f
C9137 AVDD.t6 AVSS 0.033572f
C9138 AVDD.n1282 AVSS 0.498758f
C9139 AVDD.n1283 AVSS 0.498758f
C9140 AVDD.t593 AVSS 0.089409f
C9141 AVDD.n1284 AVSS 0.55425f
C9142 AVDD.n1285 AVSS 0.49024f
C9143 AVDD.n1286 AVSS 0.021426f
C9144 AVDD.t1036 AVSS 0.021426f
C9145 AVDD.n1287 AVSS 0.021426f
C9146 AVDD.n1288 AVSS 0.49024f
C9147 AVDD.t1125 AVSS 0.089409f
C9148 AVDD.n1289 AVSS 0.55425f
C9149 AVDD.n1290 AVSS 0.49024f
C9150 AVDD.n1291 AVSS 0.021426f
C9151 AVDD.t1210 AVSS 0.033572f
C9152 AVDD.n1292 AVSS 0.515156f
C9153 AVDD.t412 AVSS 0.033572f
C9154 AVDD.t411 AVSS 0.089409f
C9155 AVDD.t1055 AVSS 0.089409f
C9156 AVDD.n1293 AVSS 0.342362f
C9157 AVDD.t549 AVSS 0.021426f
C9158 AVDD.n1294 AVSS 0.021426f
C9159 AVDD.t1173 AVSS 0.089409f
C9160 AVDD.t1174 AVSS 0.021426f
C9161 AVDD.n1295 AVSS 0.021426f
C9162 AVDD.t799 AVSS 0.089409f
C9163 AVDD.t135 AVSS 0.089409f
C9164 AVDD.n1296 AVSS 0.342362f
C9165 AVDD.t154 AVSS 0.033572f
C9166 AVDD.t800 AVSS 0.021426f
C9167 AVDD.n1297 AVSS 0.021426f
C9168 AVDD.t812 AVSS 0.089409f
C9169 AVDD.t813 AVSS 0.033572f
C9170 AVDD.t1228 AVSS 0.021426f
C9171 AVDD.n1298 AVSS 0.021426f
C9172 AVDD.t964 AVSS 0.033572f
C9173 AVDD.t963 AVSS 0.089409f
C9174 AVDD.t330 AVSS 0.089409f
C9175 AVDD.n1299 AVSS 0.342362f
C9176 AVDD.n1300 AVSS 0.021426f
C9177 AVDD.t331 AVSS 0.033572f
C9178 AVDD.n1301 AVSS 0.292092f
C9179 AVDD.n1302 AVSS 0.292092f
C9180 AVDD.t152 AVSS 0.089409f
C9181 AVDD.n1303 AVSS 0.342362f
C9182 AVDD.n1304 AVSS 0.278352f
C9183 AVDD.n1305 AVSS 0.021426f
C9184 AVDD.t137 AVSS 0.021426f
C9185 AVDD.n1306 AVSS 0.021426f
C9186 AVDD.n1307 AVSS 0.278352f
C9187 AVDD.t548 AVSS 0.089409f
C9188 AVDD.n1308 AVSS 0.342362f
C9189 AVDD.n1309 AVSS 0.278352f
C9190 AVDD.n1310 AVSS 0.021426f
C9191 AVDD.t1056 AVSS 0.033572f
C9192 AVDD.n1311 AVSS 0.301403f
C9193 AVDD.t692 AVSS 0.089409f
C9194 AVDD.t21 AVSS 0.089409f
C9195 AVDD.n1312 AVSS 0.342362f
C9196 AVDD.t693 AVSS 0.033572f
C9197 AVDD.t918 AVSS 0.021426f
C9198 AVDD.t276 AVSS 0.089409f
C9199 AVDD.t917 AVSS 0.089409f
C9200 AVDD.n1313 AVSS 0.342362f
C9201 AVDD.t553 AVSS 0.021426f
C9202 AVDD.t552 AVSS 0.089409f
C9203 AVDD.t1181 AVSS 0.089409f
C9204 AVDD.n1314 AVSS 0.342362f
C9205 AVDD.t339 AVSS 0.033572f
C9206 AVDD.t973 AVSS 0.089409f
C9207 AVDD.t337 AVSS 0.089409f
C9208 AVDD.n1315 AVSS 0.342362f
C9209 AVDD.t927 AVSS 0.089409f
C9210 AVDD.t298 AVSS 0.089409f
C9211 AVDD.n1316 AVSS 0.342362f
C9212 AVDD.t928 AVSS 0.033572f
C9213 AVDD.t568 AVSS 0.021426f
C9214 AVDD.t1193 AVSS 0.089409f
C9215 AVDD.t567 AVSS 0.089409f
C9216 AVDD.n1317 AVSS 0.218868f
C9217 AVDD.t352 AVSS 0.033572f
C9218 AVDD.t351 AVSS 0.089409f
C9219 AVDD.t993 AVSS 0.089409f
C9220 AVDD.n1318 AVSS 0.342362f
C9221 AVDD.t368 AVSS 0.089409f
C9222 AVDD.t1009 AVSS 0.089409f
C9223 AVDD.n1319 AVSS 0.342362f
C9224 AVDD.t369 AVSS 0.033572f
C9225 AVDD.t1266 AVSS 0.021426f
C9226 AVDD.t648 AVSS 0.089409f
C9227 AVDD.t1265 AVSS 0.089409f
C9228 AVDD.n1320 AVSS 0.342362f
C9229 AVDD.t1180 AVSS 0.021426f
C9230 AVDD.t1179 AVSS 0.089409f
C9231 AVDD.t559 AVSS 0.089409f
C9232 AVDD.n1321 AVSS 0.342362f
C9233 AVDD.t845 AVSS 0.033572f
C9234 AVDD.t177 AVSS 0.089409f
C9235 AVDD.t844 AVSS 0.089409f
C9236 AVDD.n1322 AVSS 0.342362f
C9237 AVDD.t179 AVSS 0.033572f
C9238 AVDD.n1323 AVSS 0.021426f
C9239 AVDD.n1324 AVSS 0.278352f
C9240 AVDD.n1325 AVSS 0.021426f
C9241 AVDD.t560 AVSS 0.021426f
C9242 AVDD.n1326 AVSS 0.021426f
C9243 AVDD.n1327 AVSS 0.278352f
C9244 AVDD.n1328 AVSS 0.021426f
C9245 AVDD.t649 AVSS 0.021426f
C9246 AVDD.n1329 AVSS 0.021426f
C9247 AVDD.n1330 AVSS 0.278352f
C9248 AVDD.n1331 AVSS 0.021426f
C9249 AVDD.t1010 AVSS 0.033572f
C9250 AVDD.n1332 AVSS 0.292092f
C9251 AVDD.n1333 AVSS 0.292092f
C9252 AVDD.t994 AVSS 0.033572f
C9253 AVDD.n1334 AVSS 0.021426f
C9254 AVDD.n1335 AVSS 0.26267f
C9255 AVDD.n1336 AVSS 0.021426f
C9256 AVDD.t1194 AVSS 0.021426f
C9257 AVDD.n1337 AVSS 0.021426f
C9258 AVDD.n1338 AVSS 0.278352f
C9259 AVDD.n1339 AVSS 0.021426f
C9260 AVDD.t299 AVSS 0.033572f
C9261 AVDD.n1340 AVSS 0.292092f
C9262 AVDD.n1341 AVSS 0.292092f
C9263 AVDD.t974 AVSS 0.033572f
C9264 AVDD.n1342 AVSS 0.021426f
C9265 AVDD.n1343 AVSS 0.278352f
C9266 AVDD.n1344 AVSS 0.021426f
C9267 AVDD.t1182 AVSS 0.021426f
C9268 AVDD.n1345 AVSS 0.021426f
C9269 AVDD.n1346 AVSS 0.278352f
C9270 AVDD.n1347 AVSS 0.021426f
C9271 AVDD.t277 AVSS 0.021426f
C9272 AVDD.n1348 AVSS 0.021426f
C9273 AVDD.n1349 AVSS 0.278352f
C9274 AVDD.n1350 AVSS 0.021426f
C9275 AVDD.t23 AVSS 0.033572f
C9276 AVDD.n1351 AVSS 0.301403f
C9277 AVDD.t391 AVSS 0.089409f
C9278 AVDD.t923 AVSS 0.089409f
C9279 AVDD.n1352 AVSS 0.70323f
C9280 AVDD.t587 AVSS 0.089409f
C9281 AVDD.t1105 AVSS 0.089409f
C9282 AVDD.n1353 AVSS 0.70323f
C9283 AVDD.t1106 AVSS 0.045717f
C9284 AVDD.t588 AVSS 0.045717f
C9285 AVDD.n1354 AVSS 1.25275f
C9286 AVDD.t1083 AVSS 0.089409f
C9287 AVDD.t349 AVSS 0.089409f
C9288 AVDD.n1355 AVSS 1.27555f
C9289 AVDD.t350 AVSS 0.045717f
C9290 AVDD.t1084 AVSS 0.045717f
C9291 AVDD.n1356 AVSS 0.720373f
C9292 AVDD.n1357 AVSS 1.08692f
C9293 AVDD.t982 AVSS 0.045717f
C9294 AVDD.t442 AVSS 0.045717f
C9295 AVDD.n1358 AVSS 0.719444f
C9296 AVDD.t441 AVSS 0.089409f
C9297 AVDD.t981 AVSS 0.089409f
C9298 AVDD.n1359 AVSS 1.27555f
C9299 AVDD.t208 AVSS 0.045717f
C9300 AVDD.t960 AVSS 0.045717f
C9301 AVDD.n1360 AVSS 1.25275f
C9302 AVDD.t959 AVSS 0.089409f
C9303 AVDD.t207 AVSS 0.089409f
C9304 AVDD.n1361 AVSS 0.70323f
C9305 AVDD.t866 AVSS 0.089409f
C9306 AVDD.t69 AVSS 0.089409f
C9307 AVDD.n1362 AVSS 0.70323f
C9308 AVDD.t71 AVSS 0.045717f
C9309 AVDD.t867 AVSS 0.045717f
C9310 AVDD.n1363 AVSS 0.872745f
C9311 AVDD.n1364 AVSS 0.378581f
C9312 AVDD.n1365 AVSS 1.19296f
C9313 AVDD.t212 AVSS 0.045717f
C9314 AVDD.t222 AVSS 0.045717f
C9315 AVDD.n1366 AVSS 0.956364f
C9316 AVDD.t221 AVSS 0.089409f
C9317 AVDD.t211 AVSS 0.089409f
C9318 AVDD.n1367 AVSS 0.70323f
C9319 AVDD.t113 AVSS 0.089409f
C9320 AVDD.t72 AVSS 0.089409f
C9321 AVDD.n1368 AVSS 0.70323f
C9322 AVDD.t73 AVSS 0.045717f
C9323 AVDD.t115 AVSS 0.045717f
C9324 AVDD.n1369 AVSS 1.25275f
C9325 AVDD.t694 AVSS 0.089409f
C9326 AVDD.t676 AVSS 0.089409f
C9327 AVDD.n1370 AVSS 1.27555f
C9328 AVDD.t677 AVSS 0.045717f
C9329 AVDD.t695 AVSS 0.045717f
C9330 AVDD.n1371 AVSS 1.2639f
C9331 AVDD.t681 AVSS 0.045717f
C9332 AVDD.t703 AVSS 0.045717f
C9333 AVDD.t702 AVSS 0.089409f
C9334 AVDD.t1178 AVSS 0.045717f
C9335 AVDD.t1192 AVSS 0.045717f
C9336 AVDD.t1191 AVSS 0.089409f
C9337 AVDD.t1069 AVSS 0.089409f
C9338 AVDD.t1059 AVSS 0.089409f
C9339 AVDD.n1372 AVSS 0.70323f
C9340 AVDD.t1177 AVSS 0.089409f
C9341 AVDD.n1373 AVSS 0.70323f
C9342 AVDD.n1374 AVSS 1.25275f
C9343 AVDD.t680 AVSS 0.089409f
C9344 AVDD.n1375 AVSS 1.27555f
C9345 AVDD.n1376 AVSS 1.26297f
C9346 AVDD.n1377 AVSS 2.38958f
C9347 AVDD.n1378 AVSS 0.515156f
C9348 AVDD.t453 AVSS 0.089409f
C9349 AVDD.n1379 AVSS 0.55425f
C9350 AVDD.n1380 AVSS 0.49024f
C9351 AVDD.n1381 AVSS 0.021426f
C9352 AVDD.t1040 AVSS 0.021426f
C9353 AVDD.n1382 AVSS 0.021426f
C9354 AVDD.n1383 AVSS 0.49024f
C9355 AVDD.t1109 AVSS 0.089409f
C9356 AVDD.n1384 AVSS 0.55425f
C9357 AVDD.n1385 AVSS 0.49024f
C9358 AVDD.n1386 AVSS 0.021426f
C9359 AVDD.t762 AVSS 0.033572f
C9360 AVDD.n1387 AVSS 0.498758f
C9361 AVDD.n1388 AVSS 0.498758f
C9362 AVDD.t157 AVSS 0.033572f
C9363 AVDD.n1389 AVSS 0.021426f
C9364 AVDD.n1390 AVSS 0.49024f
C9365 AVDD.t230 AVSS 0.089409f
C9366 AVDD.n1391 AVSS 0.33675f
C9367 AVDD.n1392 AVSS 0.24512f
C9368 AVDD.n1393 AVSS 0.374271f
C9369 AVDD.n1394 AVSS 5.09382f
C9370 AVDD.n1395 AVSS 0.378609f
C9371 AVDD.t210 AVSS 0.045717f
C9372 AVDD.t1050 AVSS 0.045717f
C9373 AVDD.n1396 AVSS 0.230382f
C9374 AVDD.t1049 AVSS 0.089409f
C9375 AVDD.t209 AVSS 0.089409f
C9376 AVDD.n1397 AVSS 0.787444f
C9377 AVDD.t730 AVSS 0.045717f
C9378 AVDD.t301 AVSS 0.045717f
C9379 AVDD.n1398 AVSS 0.764636f
C9380 AVDD.t300 AVSS 0.089409f
C9381 AVDD.t729 AVSS 0.089409f
C9382 AVDD.n1399 AVSS 0.445699f
C9383 AVDD.t166 AVSS 0.089409f
C9384 AVDD.t607 AVSS 0.089409f
C9385 AVDD.n1400 AVSS 0.445699f
C9386 AVDD.t608 AVSS 0.045717f
C9387 AVDD.t167 AVSS 0.045717f
C9388 AVDD.n1401 AVSS 0.537731f
C9389 AVDD.t685 AVSS 0.045717f
C9390 AVDD.t271 AVSS 0.045717f
C9391 AVDD.t270 AVSS 0.089409f
C9392 AVDD.t439 AVSS 0.089409f
C9393 AVDD.t894 AVSS 0.045717f
C9394 AVDD.t440 AVSS 0.045717f
C9395 AVDD.t957 AVSS 0.089409f
C9396 AVDD.t95 AVSS 0.089409f
C9397 AVDD.n1402 AVSS 0.787444f
C9398 AVDD.n1403 AVSS 0.764636f
C9399 AVDD.t893 AVSS 0.089409f
C9400 AVDD.n1404 AVSS 0.445699f
C9401 AVDD.t684 AVSS 0.089409f
C9402 AVDD.n1405 AVSS 0.445699f
C9403 AVDD.n1406 AVSS 0.587661f
C9404 AVDD.n1407 AVSS 0.712338f
C9405 AVDD.n1408 AVSS 0.375467f
C9406 AVDD.n1409 AVSS 5.56016f
C9407 AVDD.n1410 AVSS 0.375467f
C9408 AVDD.n1411 AVSS 0.712338f
C9409 AVDD.n1412 AVSS 0.537731f
C9410 AVDD.t1143 AVSS 0.089409f
C9411 AVDD.n1413 AVSS 0.445699f
C9412 AVDD.t1237 AVSS 0.089409f
C9413 AVDD.n1414 AVSS 0.445699f
C9414 AVDD.n1415 AVSS 0.764636f
C9415 AVDD.t753 AVSS 0.089409f
C9416 AVDD.n1416 AVSS 0.787444f
C9417 AVDD.n1417 AVSS 0.446192f
C9418 AVDD.n1418 AVSS 0.763137f
C9419 AVDD.n1419 AVSS 0.301403f
C9420 AVDD.t240 AVSS 0.089409f
C9421 AVDD.n1420 AVSS 0.342362f
C9422 AVDD.n1421 AVSS 0.278352f
C9423 AVDD.n1422 AVSS 0.021426f
C9424 AVDD.t661 AVSS 0.021426f
C9425 AVDD.n1423 AVSS 0.021426f
C9426 AVDD.n1424 AVSS 0.278352f
C9427 AVDD.t1033 AVSS 0.089409f
C9428 AVDD.n1425 AVSS 0.342362f
C9429 AVDD.n1426 AVSS 0.278352f
C9430 AVDD.n1427 AVSS 0.021426f
C9431 AVDD.t194 AVSS 0.033572f
C9432 AVDD.n1428 AVSS 0.292092f
C9433 AVDD.n1429 AVSS 0.292092f
C9434 AVDD.t456 AVSS 0.033572f
C9435 AVDD.n1430 AVSS 0.021426f
C9436 AVDD.n1431 AVSS 0.278352f
C9437 AVDD.t763 AVSS 0.089409f
C9438 AVDD.n1432 AVSS 0.218868f
C9439 AVDD.n1433 AVSS 0.139176f
C9440 AVDD.n1434 AVSS 0.374271f
C9441 AVDD.n1435 AVSS 5.09382f
C9442 AVDD.n1436 AVSS 0.374271f
C9443 AVDD.n1437 AVSS 0.068728f
C9444 AVDD.t870 AVSS 0.089409f
C9445 AVDD.n1438 AVSS 0.108477f
C9446 AVDD.n1439 AVSS 0.137456f
C9447 AVDD.n1440 AVSS 0.021426f
C9448 AVDD.t576 AVSS 0.033572f
C9449 AVDD.n1441 AVSS 0.144368f
C9450 AVDD.n1442 AVSS 0.144368f
C9451 AVDD.t306 AVSS 0.089409f
C9452 AVDD.n1443 AVSS 0.169461f
C9453 AVDD.n1444 AVSS 0.137456f
C9454 AVDD.n1445 AVSS 0.021426f
C9455 AVDD.t1162 AVSS 0.021426f
C9456 AVDD.n1446 AVSS 0.021426f
C9457 AVDD.n1447 AVSS 0.137456f
C9458 AVDD.t779 AVSS 0.089409f
C9459 AVDD.n1448 AVSS 0.169461f
C9460 AVDD.n1449 AVSS 0.113368f
C9461 AVDD.n1450 AVSS 0.021426f
C9462 AVDD.t345 AVSS 0.033572f
C9463 AVDD.n1451 AVSS 0.140979f
C9464 AVDD.n1452 AVSS 0.068966f
C9465 AVDD.n1453 AVSS 0.054861f
C9466 AVDD.n1454 AVSS 0.453573f
C9467 AVDD.n1455 AVSS 0.006326f
C9468 AVDD.n1456 AVSS 0.006326f
C9469 AVDD.n1457 AVSS 0.006326f
C9470 AVDD.t1506 AVSS 0.010713f
C9471 AVDD.t1541 AVSS 0.010713f
C9472 AVDD.n1458 AVSS 0.056313f
C9473 AVDD.n1459 AVSS 0.084328f
C9474 AVDD.t1357 AVSS 0.010713f
C9475 AVDD.t1326 AVSS 0.010713f
C9476 AVDD.n1460 AVSS 0.024734f
C9477 AVDD.n1461 AVSS 0.021966f
C9478 AVDD.n1462 AVSS 0.014056f
C9479 AVDD.n1463 AVSS 0.083157f
C9480 AVDD.n1464 AVSS 0.08315f
C9481 AVDD.t1347 AVSS 0.010713f
C9482 AVDD.t1336 AVSS 0.010713f
C9483 AVDD.n1465 AVSS 0.024734f
C9484 AVDD.n1466 AVSS 0.021966f
C9485 AVDD.n1467 AVSS 0.014056f
C9486 AVDD.n1468 AVSS 0.025919f
C9487 AVDD.n1469 AVSS 0.025912f
C9488 AVDD.t1514 AVSS 0.010713f
C9489 AVDD.t1343 AVSS 0.010713f
C9490 AVDD.n1470 AVSS 0.024734f
C9491 AVDD.n1471 AVSS 0.021966f
C9492 AVDD.n1472 AVSS 0.014056f
C9493 AVDD.n1473 AVSS 0.005564f
C9494 AVDD.n1474 AVSS 0.006326f
C9495 AVDD.t1632 AVSS 0.010713f
C9496 AVDD.t1376 AVSS 0.010713f
C9497 AVDD.n1475 AVSS 0.024734f
C9498 AVDD.n1476 AVSS 0.021966f
C9499 AVDD.n1477 AVSS 0.006326f
C9500 AVDD.t1372 AVSS 0.010713f
C9501 AVDD.t1606 AVSS 0.010713f
C9502 AVDD.n1478 AVSS 0.024734f
C9503 AVDD.n1479 AVSS 0.021966f
C9504 AVDD.n1480 AVSS 0.006326f
C9505 AVDD.t1553 AVSS 0.010713f
C9506 AVDD.t1315 AVSS 0.010713f
C9507 AVDD.n1481 AVSS 0.024734f
C9508 AVDD.n1482 AVSS 0.021966f
C9509 AVDD.n1483 AVSS 0.006326f
C9510 AVDD.t1621 AVSS 0.010713f
C9511 AVDD.t1368 AVSS 0.010713f
C9512 AVDD.n1484 AVSS 0.024734f
C9513 AVDD.n1485 AVSS 0.021966f
C9514 AVDD.n1486 AVSS 0.125259f
C9515 AVDD.t1354 AVSS 0.010713f
C9516 AVDD.t1608 AVSS 0.010713f
C9517 AVDD.n1487 AVSS 0.029555f
C9518 AVDD.t1522 AVSS 0.010713f
C9519 AVDD.t1615 AVSS 0.010713f
C9520 AVDD.n1488 AVSS 0.026989f
C9521 AVDD.n1489 AVSS 0.16604f
C9522 AVDD.t1504 AVSS 0.030236f
C9523 AVDD.t1623 AVSS 0.028057f
C9524 AVDD.n1490 AVSS 0.096159f
C9525 AVDD.n1491 AVSS 0.190533f
C9526 AVDD.n1492 AVSS 0.006326f
C9527 AVDD.n1493 AVSS 0.006326f
C9528 AVDD.n1494 AVSS 0.006326f
C9529 AVDD.t1501 AVSS 0.010713f
C9530 AVDD.t1511 AVSS 0.010713f
C9531 AVDD.n1495 AVSS 0.056313f
C9532 AVDD.n1496 AVSS 0.084328f
C9533 AVDD.t1311 AVSS 0.010713f
C9534 AVDD.t1319 AVSS 0.010713f
C9535 AVDD.n1497 AVSS 0.024734f
C9536 AVDD.n1498 AVSS 0.021966f
C9537 AVDD.n1499 AVSS 0.014056f
C9538 AVDD.n1500 AVSS 0.083157f
C9539 AVDD.n1501 AVSS 0.08315f
C9540 AVDD.t1544 AVSS 0.010713f
C9541 AVDD.t1498 AVSS 0.010713f
C9542 AVDD.n1502 AVSS 0.024734f
C9543 AVDD.n1503 AVSS 0.021966f
C9544 AVDD.n1504 AVSS 0.014056f
C9545 AVDD.n1505 AVSS 0.025919f
C9546 AVDD.n1506 AVSS 0.025912f
C9547 AVDD.t1508 AVSS 0.010713f
C9548 AVDD.t1332 AVSS 0.010713f
C9549 AVDD.n1507 AVSS 0.024734f
C9550 AVDD.n1508 AVSS 0.021966f
C9551 AVDD.n1509 AVSS 0.014056f
C9552 AVDD.n1510 AVSS 0.005564f
C9553 AVDD.n1511 AVSS 0.006326f
C9554 AVDD.t1349 AVSS 0.010713f
C9555 AVDD.t1359 AVSS 0.010713f
C9556 AVDD.n1512 AVSS 0.024734f
C9557 AVDD.n1513 AVSS 0.021966f
C9558 AVDD.n1514 AVSS 0.006326f
C9559 AVDD.t1535 AVSS 0.010713f
C9560 AVDD.t1543 AVSS 0.010713f
C9561 AVDD.n1515 AVSS 0.024734f
C9562 AVDD.n1516 AVSS 0.021966f
C9563 AVDD.n1517 AVSS 0.006326f
C9564 AVDD.t1512 AVSS 0.010713f
C9565 AVDD.t1335 AVSS 0.010713f
C9566 AVDD.n1518 AVSS 0.024734f
C9567 AVDD.n1519 AVSS 0.021966f
C9568 AVDD.n1520 AVSS 0.006326f
C9569 AVDD.t1610 AVSS 0.010713f
C9570 AVDD.t1546 AVSS 0.010713f
C9571 AVDD.n1521 AVSS 0.024734f
C9572 AVDD.n1522 AVSS 0.021966f
C9573 AVDD.n1523 AVSS 0.014056f
C9574 AVDD.n1524 AVSS 0.025912f
C9575 AVDD.n1525 AVSS 0.025919f
C9576 AVDD.n1526 AVSS 0.014056f
C9577 AVDD.n1527 AVSS 0.08315f
C9578 AVDD.n1528 AVSS 0.083157f
C9579 AVDD.n1529 AVSS 0.014056f
C9580 AVDD.n1530 AVSS 0.025912f
C9581 AVDD.n1531 AVSS 0.025919f
C9582 AVDD.n1532 AVSS 0.014056f
C9583 AVDD.n1533 AVSS 0.082742f
C9584 AVDD.n1534 AVSS 0.176829f
C9585 AVDD.n1535 AVSS 0.623624f
C9586 AVDD.n1536 AVSS 0.203322f
C9587 AVDD.t1308 AVSS 0.010713f
C9588 AVDD.t1634 AVSS 0.010713f
C9589 AVDD.n1537 AVSS 0.029555f
C9590 AVDD.t1317 AVSS 0.010713f
C9591 AVDD.t1560 AVSS 0.010713f
C9592 AVDD.n1538 AVSS 0.026989f
C9593 AVDD.n1539 AVSS 0.074442f
C9594 AVDD.n1540 AVSS 0.176661f
C9595 AVDD.t1377 AVSS 0.030236f
C9596 AVDD.t1346 AVSS 0.028057f
C9597 AVDD.n1541 AVSS 0.096159f
C9598 AVDD.n1542 AVSS 0.115083f
C9599 AVDD.n1543 AVSS 0.678828f
C9600 AVDD.t1331 AVSS 0.010713f
C9601 AVDD.t1638 AVSS 0.010713f
C9602 AVDD.n1544 AVSS 0.058856f
C9603 AVDD.t1532 AVSS 0.010713f
C9604 AVDD.t1345 AVSS 0.010713f
C9605 AVDD.n1545 AVSS 0.039303f
C9606 AVDD.n1546 AVSS 0.193299f
C9607 AVDD.t1523 AVSS 0.010713f
C9608 AVDD.t1355 AVSS 0.010713f
C9609 AVDD.n1547 AVSS 0.039303f
C9610 AVDD.n1548 AVSS 0.137092f
C9611 AVDD.t1337 AVSS 0.010713f
C9612 AVDD.t1518 AVSS 0.010713f
C9613 AVDD.n1549 AVSS 0.039303f
C9614 AVDD.n1550 AVSS 0.055061f
C9615 AVDD.n1551 AVSS 0.08934f
C9616 AVDD.t1314 AVSS 0.010713f
C9617 AVDD.t1618 AVSS 0.010713f
C9618 AVDD.n1552 AVSS 0.039303f
C9619 AVDD.n1553 AVSS 0.133554f
C9620 AVDD.t1550 AVSS 0.010713f
C9621 AVDD.t1362 AVSS 0.010713f
C9622 AVDD.n1554 AVSS 0.039303f
C9623 AVDD.n1555 AVSS 0.137089f
C9624 AVDD.t1509 AVSS 0.010713f
C9625 AVDD.t1559 AVSS 0.010713f
C9626 AVDD.n1556 AVSS 0.039303f
C9627 AVDD.n1557 AVSS 0.137092f
C9628 AVDD.t1305 AVSS 0.010713f
C9629 AVDD.t1542 AVSS 0.010713f
C9630 AVDD.n1558 AVSS 0.039303f
C9631 AVDD.n1559 AVSS 0.084297f
C9632 AVDD.n1560 AVSS 0.458165f
C9633 AVDD.n1561 AVSS 0.4387f
C9634 AVDD.n1562 AVSS 0.034094f
C9635 AVDD.n1563 AVSS 0.014056f
C9636 AVDD.n1564 AVSS 0.025912f
C9637 AVDD.n1565 AVSS 0.025919f
C9638 AVDD.n1566 AVSS 0.014056f
C9639 AVDD.n1567 AVSS 0.08315f
C9640 AVDD.n1568 AVSS 0.083157f
C9641 AVDD.n1569 AVSS 0.014056f
C9642 AVDD.n1570 AVSS 0.025912f
C9643 AVDD.n1571 AVSS 0.025919f
C9644 AVDD.n1572 AVSS 0.014056f
C9645 AVDD.n1573 AVSS 0.082742f
C9646 AVDD.n1574 AVSS 0.081776f
C9647 AVDD.n1575 AVSS 0.436774f
C9648 AVDD.t1622 AVSS 0.010713f
C9649 AVDD.t1534 AVSS 0.010713f
C9650 AVDD.n1576 AVSS 0.029555f
C9651 AVDD.t1612 AVSS 0.010713f
C9652 AVDD.t1526 AVSS 0.010713f
C9653 AVDD.n1577 AVSS 0.026989f
C9654 AVDD.n1578 AVSS 0.16604f
C9655 AVDD.t1348 AVSS 0.030236f
C9656 AVDD.t1562 AVSS 0.028057f
C9657 AVDD.n1579 AVSS 0.096159f
C9658 AVDD.n1580 AVSS 0.190533f
C9659 AVDD.t1373 AVSS 0.030236f
C9660 AVDD.t1363 AVSS 0.028057f
C9661 AVDD.n1581 AVSS 0.096159f
C9662 AVDD.n1582 AVSS 0.115083f
C9663 AVDD.t1505 AVSS 0.010713f
C9664 AVDD.t1556 AVSS 0.010713f
C9665 AVDD.n1583 AVSS 0.029555f
C9666 AVDD.t1495 AVSS 0.010713f
C9667 AVDD.t1551 AVSS 0.010713f
C9668 AVDD.n1584 AVSS 0.026989f
C9669 AVDD.n1585 AVSS 0.074442f
C9670 AVDD.n1586 AVSS 0.176661f
C9671 AVDD.n1587 AVSS 0.203322f
C9672 AVDD.n1588 AVSS 0.379771f
C9673 AVDD.n1589 AVSS 0.339854f
C9674 AVDD.n1590 AVSS 0.08934f
C9675 AVDD.t1513 AVSS 0.010713f
C9676 AVDD.t1547 AVSS 0.010713f
C9677 AVDD.n1591 AVSS 0.039303f
C9678 AVDD.n1592 AVSS 0.133554f
C9679 AVDD.t1325 AVSS 0.010713f
C9680 AVDD.t1629 AVSS 0.010713f
C9681 AVDD.n1593 AVSS 0.039303f
C9682 AVDD.n1594 AVSS 0.137089f
C9683 AVDD.t1350 AVSS 0.010713f
C9684 AVDD.t1338 AVSS 0.010713f
C9685 AVDD.n1595 AVSS 0.039303f
C9686 AVDD.n1596 AVSS 0.137092f
C9687 AVDD.t1502 AVSS 0.010713f
C9688 AVDD.t1320 AVSS 0.010713f
C9689 AVDD.n1597 AVSS 0.039303f
C9690 AVDD.n1598 AVSS 0.084297f
C9691 AVDD.n1599 AVSS 0.344446f
C9692 AVDD.n1600 AVSS 0.054861f
C9693 AVDD.n1601 AVSS 0.055933f
C9694 AVDD.n1602 AVSS 0.113368f
C9695 AVDD.n1603 AVSS 0.021426f
C9696 AVDD.t139 AVSS 0.033572f
C9697 AVDD.n1604 AVSS 0.140979f
C9698 AVDD.t432 AVSS 0.045717f
C9699 AVDD.t1188 AVSS 0.045717f
C9700 AVDD.n1605 AVSS 0.358025f
C9701 AVDD.n1606 AVSS 0.885941f
C9702 AVDD.n1607 AVSS 0.148966f
C9703 AVDD.t1168 AVSS 0.033572f
C9704 AVDD.t269 AVSS 0.021426f
C9705 AVDD.t286 AVSS 0.089409f
C9706 AVDD.n1608 AVSS 0.169461f
C9707 AVDD.t417 AVSS 0.089409f
C9708 AVDD.n1609 AVSS 0.169461f
C9709 AVDD.t713 AVSS 0.021426f
C9710 AVDD.t1135 AVSS 0.089409f
C9711 AVDD.n1610 AVSS 0.169461f
C9712 AVDD.t1063 AVSS 0.089409f
C9713 AVDD.n1611 AVSS 0.169461f
C9714 AVDD.t54 AVSS 0.021426f
C9715 AVDD.n1612 AVSS 0.021426f
C9716 AVDD.n1613 AVSS 0.137456f
C9717 AVDD.t52 AVSS 0.089409f
C9718 AVDD.n1614 AVSS 0.169461f
C9719 AVDD.n1615 AVSS 0.137456f
C9720 AVDD.n1616 AVSS 0.021426f
C9721 AVDD.t1064 AVSS 0.033572f
C9722 AVDD.n1617 AVSS 0.144368f
C9723 AVDD.n1618 AVSS 0.144368f
C9724 AVDD.t1136 AVSS 0.033572f
C9725 AVDD.n1619 AVSS 0.021426f
C9726 AVDD.n1620 AVSS 0.137456f
C9727 AVDD.t712 AVSS 0.089409f
C9728 AVDD.n1621 AVSS 0.108477f
C9729 AVDD.n1622 AVSS 0.068728f
C9730 AVDD.n1623 AVSS 0.129712f
C9731 AVDD.n1624 AVSS 0.021426f
C9732 AVDD.t418 AVSS 0.033572f
C9733 AVDD.n1625 AVSS 0.144368f
C9734 AVDD.n1626 AVSS 0.144368f
C9735 AVDD.t287 AVSS 0.033572f
C9736 AVDD.n1627 AVSS 0.021426f
C9737 AVDD.n1628 AVSS 0.137456f
C9738 AVDD.t268 AVSS 0.089409f
C9739 AVDD.n1629 AVSS 0.169461f
C9740 AVDD.n1630 AVSS 0.137456f
C9741 AVDD.n1631 AVSS 0.021426f
C9742 AVDD.t643 AVSS 0.021426f
C9743 AVDD.n1632 AVSS 0.021426f
C9744 AVDD.n1633 AVSS 0.117034f
C9745 AVDD.n1634 AVSS 0.06773f
C9746 AVDD.n1635 AVSS 0.519769f
C9747 AVDD.n1636 AVSS 0.006326f
C9748 AVDD.t1686 AVSS 0.027903f
C9749 AVDD.n1637 AVSS 0.038333f
C9750 AVDD.n1638 AVSS 0.006326f
C9751 AVDD.t1417 AVSS 0.010713f
C9752 AVDD.t1458 AVSS 0.010713f
C9753 AVDD.n1639 AVSS 0.026809f
C9754 AVDD.n1640 AVSS 0.027694f
C9755 AVDD.n1641 AVSS 0.006326f
C9756 AVDD.t1567 AVSS 0.027903f
C9757 AVDD.n1642 AVSS 0.038333f
C9758 AVDD.t1573 AVSS 0.010713f
C9759 AVDD.t1413 AVSS 0.010713f
C9760 AVDD.n1643 AVSS 0.092646f
C9761 AVDD.n1644 AVSS 0.199269f
C9762 AVDD.n1645 AVSS 0.014056f
C9763 AVDD.n1646 AVSS 0.054035f
C9764 AVDD.n1647 AVSS 0.006326f
C9765 AVDD.t1588 AVSS 0.027903f
C9766 AVDD.n1648 AVSS 0.038333f
C9767 AVDD.t1399 AVSS 0.010713f
C9768 AVDD.t1581 AVSS 0.010713f
C9769 AVDD.n1649 AVSS 0.092646f
C9770 AVDD.n1650 AVSS 0.199269f
C9771 AVDD.n1651 AVSS 0.014056f
C9772 AVDD.n1652 AVSS 0.054035f
C9773 AVDD.n1653 AVSS 0.283675f
C9774 AVDD.n1654 AVSS 0.006326f
C9775 AVDD.t1300 AVSS 0.027903f
C9776 AVDD.n1655 AVSS 0.038333f
C9777 AVDD.n1656 AVSS 0.006326f
C9778 AVDD.t1672 AVSS 0.010713f
C9779 AVDD.t1492 AVSS 0.010713f
C9780 AVDD.n1657 AVSS 0.026809f
C9781 AVDD.n1658 AVSS 0.027694f
C9782 AVDD.n1659 AVSS 0.149628f
C9783 AVDD.n1660 AVSS 0.014056f
C9784 AVDD.n1661 AVSS 0.025734f
C9785 AVDD.n1662 AVSS 0.025752f
C9786 AVDD.n1663 AVSS 0.014056f
C9787 AVDD.n1664 AVSS 0.128885f
C9788 AVDD.n1665 AVSS 0.715915f
C9789 AVDD.t1671 AVSS 0.010713f
C9790 AVDD.t1403 AVSS 0.010713f
C9791 AVDD.n1666 AVSS 0.03213f
C9792 AVDD.t1296 AVSS 0.010713f
C9793 AVDD.t1469 AVSS 0.010713f
C9794 AVDD.n1667 AVSS 0.024902f
C9795 AVDD.n1668 AVSS 0.073953f
C9796 AVDD.n1669 AVSS 0.06419f
C9797 AVDD.t1674 AVSS 0.010713f
C9798 AVDD.t1593 AVSS 0.010713f
C9799 AVDD.n1670 AVSS 0.03213f
C9800 AVDD.t1445 AVSS 0.010713f
C9801 AVDD.t1438 AVSS 0.010713f
C9802 AVDD.n1671 AVSS 0.024902f
C9803 AVDD.n1672 AVSS 0.073953f
C9804 AVDD.n1673 AVSS 0.115393f
C9805 AVDD.t1460 AVSS 0.010713f
C9806 AVDD.t1566 AVSS 0.010713f
C9807 AVDD.n1674 AVSS 0.03213f
C9808 AVDD.t1654 AVSS 0.010713f
C9809 AVDD.t1641 AVSS 0.010713f
C9810 AVDD.n1675 AVSS 0.024902f
C9811 AVDD.n1676 AVSS 0.073953f
C9812 AVDD.n1677 AVSS 0.115396f
C9813 AVDD.t1447 AVSS 0.010713f
C9814 AVDD.t1664 AVSS 0.010713f
C9815 AVDD.n1678 AVSS 0.03213f
C9816 AVDD.t1441 AVSS 0.010713f
C9817 AVDD.t1466 AVSS 0.010713f
C9818 AVDD.n1679 AVSS 0.024902f
C9819 AVDD.n1680 AVSS 0.073953f
C9820 AVDD.n1681 AVSS 0.113804f
C9821 AVDD.t1480 AVSS 0.010713f
C9822 AVDD.t1490 AVSS 0.010713f
C9823 AVDD.n1682 AVSS 0.03213f
C9824 AVDD.t1689 AVSS 0.010713f
C9825 AVDD.t1428 AVSS 0.010713f
C9826 AVDD.n1683 AVSS 0.024902f
C9827 AVDD.n1684 AVSS 0.103112f
C9828 AVDD.t1475 AVSS 0.010713f
C9829 AVDD.t1660 AVSS 0.010713f
C9830 AVDD.n1685 AVSS 0.03213f
C9831 AVDD.t1494 AVSS 0.010713f
C9832 AVDD.t1479 AVSS 0.010713f
C9833 AVDD.n1686 AVSS 0.024902f
C9834 AVDD.n1687 AVSS 0.073953f
C9835 AVDD.n1688 AVSS 0.148993f
C9836 AVDD.t1688 AVSS 0.010713f
C9837 AVDD.t1410 AVSS 0.010713f
C9838 AVDD.n1689 AVSS 0.03213f
C9839 AVDD.t1647 AVSS 0.010713f
C9840 AVDD.t1658 AVSS 0.010713f
C9841 AVDD.n1690 AVSS 0.024902f
C9842 AVDD.n1691 AVSS 0.073953f
C9843 AVDD.n1692 AVSS 0.115393f
C9844 AVDD.t1582 AVSS 0.010713f
C9845 AVDD.t1391 AVSS 0.010713f
C9846 AVDD.n1693 AVSS 0.03213f
C9847 AVDD.t1474 AVSS 0.010713f
C9848 AVDD.t1406 AVSS 0.010713f
C9849 AVDD.n1694 AVSS 0.024902f
C9850 AVDD.n1695 AVSS 0.073953f
C9851 AVDD.n1696 AVSS 0.030661f
C9852 AVDD.n1697 AVSS 0.0901f
C9853 AVDD.n1698 AVSS 0.632147f
C9854 AVDD.t1431 AVSS 0.010713f
C9855 AVDD.t1488 AVSS 0.010713f
C9856 AVDD.n1699 AVSS 0.042824f
C9857 AVDD.n1700 AVSS 0.156341f
C9858 AVDD.t1662 AVSS 0.04243f
C9859 AVDD.n1701 AVSS 0.202316f
C9860 AVDD.t1484 AVSS 0.082269f
C9861 AVDD.t1416 AVSS 0.010713f
C9862 AVDD.t1425 AVSS 0.010713f
C9863 AVDD.n1702 AVSS 0.042824f
C9864 AVDD.n1703 AVSS 0.289878f
C9865 AVDD.n1704 AVSS 0.203305f
C9866 AVDD.n1705 AVSS 0.453573f
C9867 AVDD.n1706 AVSS 0.406385f
C9868 AVDD.n1707 AVSS 0.197145f
C9869 AVDD.n1708 AVSS 0.149628f
C9870 AVDD.n1709 AVSS 0.014056f
C9871 AVDD.n1710 AVSS 0.025734f
C9872 AVDD.n1711 AVSS 0.025752f
C9873 AVDD.n1712 AVSS 0.014056f
C9874 AVDD.n1713 AVSS 0.081607f
C9875 AVDD.n1714 AVSS 0.447556f
C9876 AVDD.t1656 AVSS 0.010713f
C9877 AVDD.t1590 AVSS 0.010713f
C9878 AVDD.n1715 AVSS 0.03213f
C9879 AVDD.t1375 AVSS 0.010713f
C9880 AVDD.t1649 AVSS 0.010713f
C9881 AVDD.n1716 AVSS 0.024902f
C9882 AVDD.n1717 AVSS 0.103112f
C9883 AVDD.t1440 AVSS 0.010713f
C9884 AVDD.t1387 AVSS 0.010713f
C9885 AVDD.n1718 AVSS 0.03213f
C9886 AVDD.t1432 AVSS 0.010713f
C9887 AVDD.t1489 AVSS 0.010713f
C9888 AVDD.n1719 AVSS 0.024902f
C9889 AVDD.n1720 AVSS 0.073953f
C9890 AVDD.n1721 AVSS 0.148993f
C9891 AVDD.t1450 AVSS 0.010713f
C9892 AVDD.t1569 AVSS 0.010713f
C9893 AVDD.n1722 AVSS 0.03213f
C9894 AVDD.t1476 AVSS 0.010713f
C9895 AVDD.t1690 AVSS 0.010713f
C9896 AVDD.n1723 AVSS 0.024902f
C9897 AVDD.n1724 AVSS 0.073953f
C9898 AVDD.n1725 AVSS 0.115393f
C9899 AVDD.t1463 AVSS 0.010713f
C9900 AVDD.t1680 AVSS 0.010713f
C9901 AVDD.n1726 AVSS 0.03213f
C9902 AVDD.t1293 AVSS 0.010713f
C9903 AVDD.t1592 AVSS 0.010713f
C9904 AVDD.n1727 AVSS 0.024902f
C9905 AVDD.n1728 AVSS 0.073953f
C9906 AVDD.n1729 AVSS 0.030661f
C9907 AVDD.n1730 AVSS 0.0901f
C9908 AVDD.t1424 AVSS 0.010713f
C9909 AVDD.t1397 AVSS 0.010713f
C9910 AVDD.n1731 AVSS 0.03213f
C9911 AVDD.t1437 AVSS 0.010713f
C9912 AVDD.t1383 AVSS 0.010713f
C9913 AVDD.n1732 AVSS 0.024902f
C9914 AVDD.n1733 AVSS 0.073953f
C9915 AVDD.n1734 AVSS 0.113804f
C9916 AVDD.t1429 AVSS 0.010713f
C9917 AVDD.t1485 AVSS 0.010713f
C9918 AVDD.n1735 AVSS 0.03213f
C9919 AVDD.t1405 AVSS 0.010713f
C9920 AVDD.t1451 AVSS 0.010713f
C9921 AVDD.n1736 AVSS 0.024902f
C9922 AVDD.n1737 AVSS 0.073953f
C9923 AVDD.n1738 AVSS 0.115396f
C9924 AVDD.t1473 AVSS 0.010713f
C9925 AVDD.t1468 AVSS 0.010713f
C9926 AVDD.n1739 AVSS 0.03213f
C9927 AVDD.t1462 AVSS 0.010713f
C9928 AVDD.t1303 AVSS 0.010713f
C9929 AVDD.n1740 AVSS 0.024902f
C9930 AVDD.n1741 AVSS 0.073953f
C9931 AVDD.n1742 AVSS 0.115393f
C9932 AVDD.t1404 AVSS 0.010713f
C9933 AVDD.t1563 AVSS 0.010713f
C9934 AVDD.n1743 AVSS 0.03213f
C9935 AVDD.t1393 AVSS 0.010713f
C9936 AVDD.t1682 AVSS 0.010713f
C9937 AVDD.n1744 AVSS 0.024902f
C9938 AVDD.n1745 AVSS 0.073953f
C9939 AVDD.n1746 AVSS 0.06419f
C9940 AVDD.n1747 AVSS 0.413506f
C9941 AVDD.n1748 AVSS 0.434267f
C9942 AVDD.t1578 AVSS 0.010713f
C9943 AVDD.t1586 AVSS 0.010713f
C9944 AVDD.n1749 AVSS 0.042824f
C9945 AVDD.n1750 AVSS 0.156341f
C9946 AVDD.t1394 AVSS 0.04243f
C9947 AVDD.n1751 AVSS 0.202316f
C9948 AVDD.t1583 AVSS 0.082269f
C9949 AVDD.t1667 AVSS 0.010713f
C9950 AVDD.t1289 AVSS 0.010713f
C9951 AVDD.n1752 AVSS 0.042824f
C9952 AVDD.n1753 AVSS 0.289878f
C9953 AVDD.n1754 AVSS 0.203305f
C9954 AVDD.n1755 AVSS 0.368072f
C9955 AVDD.n1756 AVSS 0.06773f
C9956 AVDD.n1757 AVSS 0.117034f
C9957 AVDD.n1758 AVSS 0.021426f
C9958 AVDD.t738 AVSS 0.021426f
C9959 AVDD.n1759 AVSS 0.021426f
C9960 AVDD.n1760 AVSS 0.137456f
C9961 AVDD.t145 AVSS 0.089409f
C9962 AVDD.n1761 AVSS 0.169461f
C9963 AVDD.n1762 AVSS 0.137456f
C9964 AVDD.n1763 AVSS 0.021426f
C9965 AVDD.t586 AVSS 0.033572f
C9966 AVDD.n1764 AVSS 0.144368f
C9967 AVDD.n1765 AVSS 0.144368f
C9968 AVDD.t343 AVSS 0.033572f
C9969 AVDD.n1766 AVSS 0.021426f
C9970 AVDD.n1767 AVSS 0.129712f
C9971 AVDD.n1768 AVSS 0.068728f
C9972 AVDD.t304 AVSS 0.089409f
C9973 AVDD.n1769 AVSS 0.108477f
C9974 AVDD.n1770 AVSS 0.137456f
C9975 AVDD.n1771 AVSS 0.021426f
C9976 AVDD.t732 AVSS 0.033572f
C9977 AVDD.n1772 AVSS 0.144368f
C9978 AVDD.n1773 AVSS 0.144368f
C9979 AVDD.t995 AVSS 0.089409f
C9980 AVDD.n1774 AVSS 0.169461f
C9981 AVDD.n1775 AVSS 0.137456f
C9982 AVDD.n1776 AVSS 0.021426f
C9983 AVDD.t1248 AVSS 0.021426f
C9984 AVDD.n1777 AVSS 0.021426f
C9985 AVDD.n1778 AVSS 0.137456f
C9986 AVDD.t868 AVSS 0.089409f
C9987 AVDD.n1779 AVSS 0.169461f
C9988 AVDD.n1780 AVSS 0.113368f
C9989 AVDD.n1781 AVSS 0.021426f
C9990 AVDD.t819 AVSS 0.033572f
C9991 AVDD.n1782 AVSS 0.174655f
C9992 AVDD.n1783 AVSS 0.068966f
C9993 AVDD.n1784 AVSS 0.054861f
C9994 AVDD.n1785 AVSS 0.458165f
C9995 AVDD.n1786 AVSS 0.006326f
C9996 AVDD.n1787 AVSS 0.006326f
C9997 AVDD.n1788 AVSS 0.006326f
C9998 AVDD.n1789 AVSS 0.006326f
C9999 AVDD.n1790 AVSS 0.006326f
C10000 AVDD.n1791 AVSS 0.006326f
C10001 AVDD.n1792 AVSS 0.006326f
C10002 AVDD.t1452 AVSS 0.010713f
C10003 AVDD.t1643 AVSS 0.010713f
C10004 AVDD.n1793 AVSS 0.056313f
C10005 AVDD.n1794 AVSS 0.084328f
C10006 AVDD.t1659 AVSS 0.010713f
C10007 AVDD.t1577 AVSS 0.010713f
C10008 AVDD.n1795 AVSS 0.024734f
C10009 AVDD.n1796 AVSS 0.021966f
C10010 AVDD.n1797 AVSS 0.014056f
C10011 AVDD.n1798 AVSS 0.083157f
C10012 AVDD.n1799 AVSS 0.08315f
C10013 AVDD.t1487 AVSS 0.010713f
C10014 AVDD.t1301 AVSS 0.010713f
C10015 AVDD.n1800 AVSS 0.024734f
C10016 AVDD.n1801 AVSS 0.021966f
C10017 AVDD.n1802 AVSS 0.014056f
C10018 AVDD.n1803 AVSS 0.025919f
C10019 AVDD.n1804 AVSS 0.025912f
C10020 AVDD.t1398 AVSS 0.010713f
C10021 AVDD.t1443 AVSS 0.010713f
C10022 AVDD.n1805 AVSS 0.024734f
C10023 AVDD.n1806 AVSS 0.021966f
C10024 AVDD.n1807 AVSS 0.014056f
C10025 AVDD.n1808 AVSS 0.005564f
C10026 AVDD.n1809 AVSS 0.006326f
C10027 AVDD.n1810 AVSS 0.006326f
C10028 AVDD.n1811 AVSS 0.006326f
C10029 AVDD.t1472 AVSS 0.010713f
C10030 AVDD.t1454 AVSS 0.010713f
C10031 AVDD.n1812 AVSS 0.056313f
C10032 AVDD.n1813 AVSS 0.084328f
C10033 AVDD.t1483 AVSS 0.010713f
C10034 AVDD.t1645 AVSS 0.010713f
C10035 AVDD.n1814 AVSS 0.024734f
C10036 AVDD.n1815 AVSS 0.021966f
C10037 AVDD.n1816 AVSS 0.014056f
C10038 AVDD.n1817 AVSS 0.083157f
C10039 AVDD.n1818 AVSS 0.08315f
C10040 AVDD.t1679 AVSS 0.010713f
C10041 AVDD.t1589 AVSS 0.010713f
C10042 AVDD.n1819 AVSS 0.024734f
C10043 AVDD.n1820 AVSS 0.021966f
C10044 AVDD.n1821 AVSS 0.014056f
C10045 AVDD.n1822 AVSS 0.025919f
C10046 AVDD.n1823 AVSS 0.025912f
C10047 AVDD.t1477 AVSS 0.010713f
C10048 AVDD.t1448 AVSS 0.010713f
C10049 AVDD.n1824 AVSS 0.024734f
C10050 AVDD.n1825 AVSS 0.021966f
C10051 AVDD.n1826 AVSS 0.014056f
C10052 AVDD.n1827 AVSS 0.005564f
C10053 AVDD.n1828 AVSS 0.176829f
C10054 AVDD.t1421 AVSS 0.010713f
C10055 AVDD.t1395 AVSS 0.010713f
C10056 AVDD.n1829 AVSS 0.029555f
C10057 AVDD.t1665 AVSS 0.010713f
C10058 AVDD.t1657 AVSS 0.010713f
C10059 AVDD.n1830 AVSS 0.026989f
C10060 AVDD.n1831 AVSS 0.16604f
C10061 AVDD.t1292 AVSS 0.030236f
C10062 AVDD.t1453 AVSS 0.028057f
C10063 AVDD.n1832 AVSS 0.096159f
C10064 AVDD.n1833 AVSS 0.190533f
C10065 AVDD.n1834 AVSS 0.006326f
C10066 AVDD.n1835 AVSS 0.006326f
C10067 AVDD.n1836 AVSS 0.006326f
C10068 AVDD.n1837 AVSS 0.006326f
C10069 AVDD.n1838 AVSS 0.082742f
C10070 AVDD.t1456 AVSS 0.010713f
C10071 AVDD.t1435 AVSS 0.010713f
C10072 AVDD.n1839 AVSS 0.024734f
C10073 AVDD.n1840 AVSS 0.021966f
C10074 AVDD.n1841 AVSS 0.014056f
C10075 AVDD.n1842 AVSS 0.025919f
C10076 AVDD.n1843 AVSS 0.025912f
C10077 AVDD.t1596 AVSS 0.010713f
C10078 AVDD.t1286 AVSS 0.010713f
C10079 AVDD.n1844 AVSS 0.024734f
C10080 AVDD.n1845 AVSS 0.021966f
C10081 AVDD.n1846 AVSS 0.014056f
C10082 AVDD.n1847 AVSS 0.083157f
C10083 AVDD.n1848 AVSS 0.08315f
C10084 AVDD.t1400 AVSS 0.010713f
C10085 AVDD.t1388 AVSS 0.010713f
C10086 AVDD.n1849 AVSS 0.024734f
C10087 AVDD.n1850 AVSS 0.021966f
C10088 AVDD.n1851 AVSS 0.014056f
C10089 AVDD.n1852 AVSS 0.025919f
C10090 AVDD.n1853 AVSS 0.025912f
C10091 AVDD.t1571 AVSS 0.010713f
C10092 AVDD.t1419 AVSS 0.010713f
C10093 AVDD.n1854 AVSS 0.024734f
C10094 AVDD.n1855 AVSS 0.021966f
C10095 AVDD.n1856 AVSS 0.014056f
C10096 AVDD.n1857 AVSS 0.125259f
C10097 AVDD.n1858 AVSS 0.678827f
C10098 AVDD.t1392 AVSS 0.030236f
C10099 AVDD.t1422 AVSS 0.028057f
C10100 AVDD.n1859 AVSS 0.096159f
C10101 AVDD.n1860 AVSS 0.115083f
C10102 AVDD.t1652 AVSS 0.010713f
C10103 AVDD.t1584 AVSS 0.010713f
C10104 AVDD.n1861 AVSS 0.029555f
C10105 AVDD.t1374 AVSS 0.010713f
C10106 AVDD.t1493 AVSS 0.010713f
C10107 AVDD.n1862 AVSS 0.026989f
C10108 AVDD.n1863 AVSS 0.074442f
C10109 AVDD.n1864 AVSS 0.176661f
C10110 AVDD.n1865 AVSS 0.203322f
C10111 AVDD.n1866 AVSS 0.623624f
C10112 AVDD.t1579 AVSS 0.010713f
C10113 AVDD.t1385 AVSS 0.010713f
C10114 AVDD.n1867 AVSS 0.058856f
C10115 AVDD.t1648 AVSS 0.010713f
C10116 AVDD.t1644 AVSS 0.010713f
C10117 AVDD.n1868 AVSS 0.039303f
C10118 AVDD.n1869 AVSS 0.193299f
C10119 AVDD.t1668 AVSS 0.010713f
C10120 AVDD.t1681 AVSS 0.010713f
C10121 AVDD.n1870 AVSS 0.039303f
C10122 AVDD.n1871 AVSS 0.137092f
C10123 AVDD.t1464 AVSS 0.010713f
C10124 AVDD.t1570 AVSS 0.010713f
C10125 AVDD.n1872 AVSS 0.039303f
C10126 AVDD.n1873 AVSS 0.055061f
C10127 AVDD.t1442 AVSS 0.010713f
C10128 AVDD.t1449 AVSS 0.010713f
C10129 AVDD.n1874 AVSS 0.039303f
C10130 AVDD.n1875 AVSS 0.084297f
C10131 AVDD.t1299 AVSS 0.010713f
C10132 AVDD.t1564 AVSS 0.010713f
C10133 AVDD.n1876 AVSS 0.039303f
C10134 AVDD.n1877 AVSS 0.137092f
C10135 AVDD.t1591 AVSS 0.010713f
C10136 AVDD.t1396 AVSS 0.010713f
C10137 AVDD.n1878 AVSS 0.039303f
C10138 AVDD.n1879 AVSS 0.137089f
C10139 AVDD.t1423 AVSS 0.010713f
C10140 AVDD.t1482 AVSS 0.010713f
C10141 AVDD.n1880 AVSS 0.039303f
C10142 AVDD.n1881 AVSS 0.133554f
C10143 AVDD.n1882 AVSS 0.08934f
C10144 AVDD.n1883 AVSS 0.453573f
C10145 AVDD.n1884 AVSS 0.436774f
C10146 AVDD.n1885 AVSS 0.081776f
C10147 AVDD.n1886 AVSS 0.082742f
C10148 AVDD.t1572 AVSS 0.010713f
C10149 AVDD.t1439 AVSS 0.010713f
C10150 AVDD.n1887 AVSS 0.024734f
C10151 AVDD.n1888 AVSS 0.021966f
C10152 AVDD.n1889 AVSS 0.014056f
C10153 AVDD.n1890 AVSS 0.025919f
C10154 AVDD.n1891 AVSS 0.025912f
C10155 AVDD.t1669 AVSS 0.010713f
C10156 AVDD.t1655 AVSS 0.010713f
C10157 AVDD.n1892 AVSS 0.024734f
C10158 AVDD.n1893 AVSS 0.021966f
C10159 AVDD.n1894 AVSS 0.014056f
C10160 AVDD.n1895 AVSS 0.083157f
C10161 AVDD.n1896 AVSS 0.08315f
C10162 AVDD.t1389 AVSS 0.010713f
C10163 AVDD.t1470 AVSS 0.010713f
C10164 AVDD.n1897 AVSS 0.024734f
C10165 AVDD.n1898 AVSS 0.021966f
C10166 AVDD.n1899 AVSS 0.014056f
C10167 AVDD.n1900 AVSS 0.025919f
C10168 AVDD.n1901 AVSS 0.025912f
C10169 AVDD.t1409 AVSS 0.010713f
C10170 AVDD.t1430 AVSS 0.010713f
C10171 AVDD.n1902 AVSS 0.024734f
C10172 AVDD.n1903 AVSS 0.021966f
C10173 AVDD.n1904 AVSS 0.014056f
C10174 AVDD.n1905 AVSS 0.034094f
C10175 AVDD.n1906 AVSS 0.4387f
C10176 AVDD.t1670 AVSS 0.010713f
C10177 AVDD.t1684 AVSS 0.010713f
C10178 AVDD.n1907 AVSS 0.029555f
C10179 AVDD.t1661 AVSS 0.010713f
C10180 AVDD.t1675 AVSS 0.010713f
C10181 AVDD.n1908 AVSS 0.026989f
C10182 AVDD.n1909 AVSS 0.16604f
C10183 AVDD.t1408 AVSS 0.030236f
C10184 AVDD.t1401 AVSS 0.028057f
C10185 AVDD.n1910 AVSS 0.096159f
C10186 AVDD.n1911 AVSS 0.190533f
C10187 AVDD.n1912 AVSS 0.203322f
C10188 AVDD.t1459 AVSS 0.010713f
C10189 AVDD.t1465 AVSS 0.010713f
C10190 AVDD.n1913 AVSS 0.029555f
C10191 AVDD.t1288 AVSS 0.010713f
C10192 AVDD.t1295 AVSS 0.010713f
C10193 AVDD.n1914 AVSS 0.026989f
C10194 AVDD.n1915 AVSS 0.074442f
C10195 AVDD.n1916 AVSS 0.176661f
C10196 AVDD.t1683 AVSS 0.030236f
C10197 AVDD.t1594 AVSS 0.028057f
C10198 AVDD.n1917 AVSS 0.096159f
C10199 AVDD.n1918 AVSS 0.115083f
C10200 AVDD.n1919 AVSS 0.429161f
C10201 AVDD.n1920 AVSS 0.344446f
C10202 AVDD.t1420 AVSS 0.010713f
C10203 AVDD.t1642 AVSS 0.010713f
C10204 AVDD.n1921 AVSS 0.039303f
C10205 AVDD.n1922 AVSS 0.084297f
C10206 AVDD.t1411 AVSS 0.010713f
C10207 AVDD.t1478 AVSS 0.010713f
C10208 AVDD.n1923 AVSS 0.039303f
C10209 AVDD.n1924 AVSS 0.137092f
C10210 AVDD.t1467 AVSS 0.010713f
C10211 AVDD.t1687 AVSS 0.010713f
C10212 AVDD.n1925 AVSS 0.039303f
C10213 AVDD.n1926 AVSS 0.137089f
C10214 AVDD.t1673 AVSS 0.010713f
C10215 AVDD.t1580 AVSS 0.010713f
C10216 AVDD.n1927 AVSS 0.039303f
C10217 AVDD.n1928 AVSS 0.133554f
C10218 AVDD.n1929 AVSS 0.08934f
C10219 AVDD.n1930 AVSS 0.339854f
C10220 AVDD.n1931 AVSS 0.054861f
C10221 AVDD.n1932 AVSS 0.055933f
C10222 AVDD.n1933 AVSS 0.113368f
C10223 AVDD.n1934 AVSS 0.021426f
C10224 AVDD.t1208 AVSS 0.033572f
C10225 AVDD.n1935 AVSS 0.140979f
C10226 AVDD.n1936 AVSS 0.585364f
C10227 AVDD.t47 AVSS 0.045717f
C10228 AVDD.t169 AVSS 0.045717f
C10229 AVDD.n1937 AVSS 0.230382f
C10230 AVDD.t168 AVSS 0.089409f
C10231 AVDD.t46 AVSS 0.089409f
C10232 AVDD.n1938 AVSS 0.787444f
C10233 AVDD.t584 AVSS 0.045717f
C10234 AVDD.t691 AVSS 0.045717f
C10235 AVDD.n1939 AVSS 0.764636f
C10236 AVDD.t690 AVSS 0.089409f
C10237 AVDD.t583 AVSS 0.089409f
C10238 AVDD.n1940 AVSS 0.445699f
C10239 AVDD.t577 AVSS 0.089409f
C10240 AVDD.t451 AVSS 0.089409f
C10241 AVDD.n1941 AVSS 0.445699f
C10242 AVDD.t452 AVSS 0.045717f
C10243 AVDD.t578 AVSS 0.045717f
C10244 AVDD.n1942 AVSS 0.537731f
C10245 AVDD.n1943 AVSS 0.378581f
C10246 AVDD.t551 AVSS 0.045717f
C10247 AVDD.t651 AVSS 0.045717f
C10248 AVDD.t650 AVSS 0.089409f
C10249 AVDD.t862 AVSS 0.089409f
C10250 AVDD.t752 AVSS 0.045717f
C10251 AVDD.t863 AVSS 0.045717f
C10252 AVDD.t48 AVSS 0.089409f
C10253 AVDD.t1235 AVSS 0.089409f
C10254 AVDD.n1944 AVSS 0.787444f
C10255 AVDD.n1945 AVSS 0.764636f
C10256 AVDD.t751 AVSS 0.089409f
C10257 AVDD.n1946 AVSS 0.445699f
C10258 AVDD.t550 AVSS 0.089409f
C10259 AVDD.n1947 AVSS 0.445699f
C10260 AVDD.n1948 AVSS 0.587661f
C10261 AVDD.n1949 AVSS 0.712338f
C10262 AVDD.n1950 AVSS 0.375467f
C10263 AVDD.n1951 AVSS 5.56016f
C10264 AVDD.n1952 AVSS 0.375467f
C10265 AVDD.n1953 AVSS 0.712338f
C10266 AVDD.n1954 AVSS 0.537731f
C10267 AVDD.t999 AVSS 0.089409f
C10268 AVDD.n1955 AVSS 0.445699f
C10269 AVDD.t1099 AVSS 0.089409f
C10270 AVDD.n1956 AVSS 0.445699f
C10271 AVDD.n1957 AVSS 0.764636f
C10272 AVDD.t605 AVSS 0.089409f
C10273 AVDD.n1958 AVSS 0.787444f
C10274 AVDD.n1959 AVSS 0.446192f
C10275 AVDD.n1960 AVSS 0.763137f
C10276 AVDD.n1961 AVSS 0.301403f
C10277 AVDD.t1111 AVSS 0.089409f
C10278 AVDD.n1962 AVSS 0.342362f
C10279 AVDD.n1963 AVSS 0.278352f
C10280 AVDD.n1964 AVSS 0.021426f
C10281 AVDD.t853 AVSS 0.021426f
C10282 AVDD.n1965 AVSS 0.021426f
C10283 AVDD.n1966 AVSS 0.278352f
C10284 AVDD.t1241 AVSS 0.089409f
C10285 AVDD.n1967 AVSS 0.342362f
C10286 AVDD.n1968 AVSS 0.278352f
C10287 AVDD.n1969 AVSS 0.021426f
C10288 AVDD.t988 AVSS 0.033572f
C10289 AVDD.n1970 AVSS 0.292092f
C10290 AVDD.n1971 AVSS 0.292092f
C10291 AVDD.t1024 AVSS 0.033572f
C10292 AVDD.n1972 AVSS 0.021426f
C10293 AVDD.n1973 AVSS 0.278352f
C10294 AVDD.t609 AVSS 0.089409f
C10295 AVDD.n1974 AVSS 0.218868f
C10296 AVDD.n1975 AVSS 0.139176f
C10297 AVDD.n1976 AVSS 0.374271f
C10298 AVDD.n1977 AVSS 5.09382f
C10299 AVDD.n1978 AVSS 0.378609f
C10300 AVDD.n1979 AVSS 0.07081f
C10301 AVDD.n1980 AVSS 0.133642f
C10302 AVDD.n1981 AVSS 0.021426f
C10303 AVDD.t356 AVSS 0.033572f
C10304 AVDD.n1982 AVSS 0.148431f
C10305 AVDD.n1983 AVSS 0.148431f
C10306 AVDD.t183 AVSS 0.089409f
C10307 AVDD.n1984 AVSS 0.173626f
C10308 AVDD.n1985 AVSS 0.141621f
C10309 AVDD.n1986 AVSS 0.021426f
C10310 AVDD.t171 AVSS 0.021426f
C10311 AVDD.n1987 AVSS 0.021426f
C10312 AVDD.n1988 AVSS 0.141621f
C10313 AVDD.t571 AVSS 0.089409f
C10314 AVDD.n1989 AVSS 0.173626f
C10315 AVDD.n1990 AVSS 0.141621f
C10316 AVDD.n1991 AVSS 0.021426f
C10317 AVDD.t1074 AVSS 0.033572f
C10318 AVDD.n1992 AVSS 0.153168f
C10319 AVDD.n1993 AVSS 0.921769f
C10320 AVDD.n1994 AVSS 0.369174f
C10321 AVDD.t370 AVSS 0.089409f
C10322 AVDD.n1995 AVSS 1.27555f
C10323 AVDD.n1996 AVSS 1.25275f
C10324 AVDD.t889 AVSS 0.089409f
C10325 AVDD.n1997 AVSS 0.70323f
C10326 AVDD.t781 AVSS 0.089409f
C10327 AVDD.n1998 AVSS 0.70323f
C10328 AVDD.n1999 AVSS 0.956364f
C10329 AVDD.n2000 AVSS 1.19296f
C10330 AVDD.n2001 AVSS 0.872745f
C10331 AVDD.t793 AVSS 0.089409f
C10332 AVDD.n2002 AVSS 0.70323f
C10333 AVDD.t668 AVSS 0.089409f
C10334 AVDD.n2003 AVSS 0.70323f
C10335 AVDD.n2004 AVSS 1.25275f
C10336 AVDD.t1225 AVSS 0.089409f
C10337 AVDD.n2005 AVSS 1.27555f
C10338 AVDD.n2006 AVSS 0.719444f
C10339 AVDD.n2007 AVSS 1.08692f
C10340 AVDD.n2008 AVSS 0.720373f
C10341 AVDD.t848 AVSS 0.089409f
C10342 AVDD.n2009 AVSS 1.27555f
C10343 AVDD.n2010 AVSS 1.25275f
C10344 AVDD.t759 AVSS 0.089409f
C10345 AVDD.n2011 AVSS 0.70323f
C10346 AVDD.t1065 AVSS 0.089409f
C10347 AVDD.n2012 AVSS 0.70323f
C10348 AVDD.n2013 AVSS 0.956364f
C10349 AVDD.n2014 AVSS 1.19296f
C10350 AVDD.n2015 AVSS 0.375467f
C10351 AVDD.n2016 AVSS 16.0886f
C10352 AVDD.n2017 AVSS 0.375467f
C10353 AVDD.n2018 AVSS 1.19296f
C10354 AVDD.n2019 AVSS 0.872745f
C10355 AVDD.t854 AVSS 0.089409f
C10356 AVDD.n2020 AVSS 0.70323f
C10357 AVDD.t953 AVSS 0.089409f
C10358 AVDD.n2021 AVSS 0.70323f
C10359 AVDD.n2022 AVSS 0.852305f
.ends

