* NGSPICE file created from CM_nfets.ext - technology: gf180mcuD

.subckt CM_nfets VSS OUT1 OUT2 IN
X0 a_n522_n1809# IN a_n1082_n1809# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1 a_352_1779# IN a_n170_882# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2 a_2346_n15# IN a_1786_882# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3 a_1786_n15# IN a_1264_n1809# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5 a_1786_n3603# IN a_1264_n3603# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6 a_912_n4500# IN a_352_n4500# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X7 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X8 a_n1082_n1809# IN a_n1604_n2706# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X9 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X10 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X11 a_352_n2706# IN a_n170_n3603# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X12 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X13 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X14 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X15 a_2346_1779# IN a_1786_2676# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X16 a_n522_882# IN a_n1082_1779# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X17 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X18 a_n1082_1779# IN a_n1604_1779# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X19 a_1786_1779# IN a_1264_882# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X20 a_912_882# IN a_352_882# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X21 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X22 a_2346_n2706# IN a_1786_n2706# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X23 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X24 a_1786_n4500# IN a_n522_n4500# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X25 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X26 a_912_1779# IN a_352_1779# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X27 a_2346_n15# IN a_1786_n15# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X28 a_n522_n3603# IN a_n1082_n2706# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X29 a_352_2676# IN a_n522_n912# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X30 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X31 IN IN VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X32 a_n1082_n2706# IN a_n1604_n2706# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X33 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X34 a_352_n3603# IN a_n170_n3603# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X35 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X36 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X37 OUT1 IN a_n1082_2676# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X38 IN IN VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X39 a_1786_2676# IN VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X40 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X41 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X42 a_2346_n4500# IN a_1786_n3603# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X43 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X44 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X45 a_n1082_2676# IN a_n1604_1779# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X46 a_1786_n1809# IN a_1264_n1809# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X47 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X48 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X49 a_912_1779# IN a_352_2676# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X50 a_n1082_882# IN a_n1604_n15# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X51 a_n522_n3603# IN a_n1082_n3603# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X52 a_352_n4500# IN VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X53 a_912_n2706# IN a_1786_n912# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X54 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X55 a_912_n2706# IN a_352_n2706# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X56 a_n1082_n3603# IN a_n1604_n4500# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X57 a_n522_882# IN a_n1082_882# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X58 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X59 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X60 a_2346_n4500# IN a_1786_n4500# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X61 VSS IN IN VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X62 a_352_882# IN a_n170_882# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X63 a_n522_n4500# IN a_n1082_n4500# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X64 a_n1082_n15# IN a_n1604_n15# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X65 a_1786_n2706# IN a_1264_n3603# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X66 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X67 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X68 a_n1082_n4500# IN a_n1604_n4500# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X69 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X70 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X71 a_1786_882# IN a_1264_882# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X72 a_n522_n912# IN a_n1082_n912# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X73 a_1786_n912# IN a_912_882# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X74 VSS IN IN VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X75 a_n522_n1809# IN a_n1082_n15# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X76 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X77 a_n1082_n912# IN OUT2 VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X78 a_912_n4500# IN a_352_n3603# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X79 a_2346_1779# IN a_1786_1779# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X80 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X81 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X82 IN IN VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X83 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X84 VSS IN IN VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X85 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X86 a_2346_n2706# IN a_1786_n1809# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X87 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
.ends

