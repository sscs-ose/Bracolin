* Extracted by KLayout with GF180MCU LVS runset on : 29/11/2023 19:35

.SUBCKT FC_pfets D1 S1 G1 G2 D2 S2 B
M$1 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$4 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$5 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$6 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$7 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$8 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$9 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$10 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$11 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$12 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$13 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$14 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$15 S1 G1 D1 B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$16 D1 G1 S1 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$17 S1 G1 D1 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$18 D1 G1 S1 B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$19 S2 G2 D2 B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$20 D2 G2 S2 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$21 S2 G2 D2 B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$22 S1 G1 D1 B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$23 D1 G1 S1 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$24 S1 G1 D1 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$25 D1 G1 S1 B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$26 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$27 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$28 S2 G2 D2 B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$29 D2 G2 S2 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$30 S2 G2 D2 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$31 D2 G2 S2 B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$32 D1 G1 S1 B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$33 S1 G1 D1 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$34 D1 G1 S1 B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$35 S2 G2 D2 B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$36 D2 G2 S2 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$37 S2 G2 D2 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$38 D2 G2 S2 B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$39 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$40 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$41 S2 G2 D2 B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$42 D2 G2 S2 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$43 S2 G2 D2 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$44 D2 G2 S2 B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$45 D1 G1 S1 B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$46 S1 G1 D1 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$47 D1 G1 S1 B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$48 S2 G2 D2 B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$49 D2 G2 S2 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$50 S2 G2 D2 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$51 D2 G2 S2 B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$52 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$53 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$54 S1 G1 D1 B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$55 D1 G1 S1 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$56 S1 G1 D1 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$57 D1 G1 S1 B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$58 D2 G2 S2 B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$59 S2 G2 D2 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$60 D2 G2 S2 B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$61 S1 G1 D1 B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$62 D1 G1 S1 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$63 S1 G1 D1 B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$64 D1 G1 S1 B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$65 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$66 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$67 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$68 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$69 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$70 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$71 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$72 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$73 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$74 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$75 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$76 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$77 B B B B pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$78 B B B B pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
.ENDS FC_pfets
