* Extracted by KLayout with GF180MCU LVS runset on : 08/04/2024 20:27

.SUBCKT UndervoltageProtection GND PowerGate vdd vfb vref iref
M$1 \$31 vfb \$5 vdd pfet_03v3 L=2U W=2U AS=1.3P AD=0.52P PS=5.3U PD=2.52U
M$2 \$5 vfb \$31 vdd pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$3 \$31 vfb \$5 vdd pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$4 \$5 vfb \$31 vdd pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$5 \$31 vfb \$5 vdd pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$6 \$5 vfb \$31 vdd pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$7 \$31 vfb \$5 vdd pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$8 \$5 vfb \$31 vdd pfet_03v3 L=2U W=2U AS=0.52P AD=1.3P PS=2.52U PD=5.3U
M$9 \$31 vref GND vdd pfet_03v3 L=2U W=2U AS=1.3P AD=0.52P PS=5.3U PD=2.52U
M$10 GND vref \$31 vdd pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$11 \$31 vref GND vdd pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$12 GND vref \$31 vdd pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$13 \$31 vref GND vdd pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$14 GND vref \$31 vdd pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$15 \$31 vref GND vdd pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$16 GND vref \$31 vdd pfet_03v3 L=2U W=2U AS=0.52P AD=1.3P PS=2.52U PD=5.3U
M$17 vdd iref \$4 vdd pfet_03v3 L=2U W=2U AS=1.3P AD=0.52P PS=5.3U PD=2.52U
M$18 \$4 iref vdd vdd pfet_03v3 L=2U W=2U AS=0.52P AD=1.3P PS=2.52U PD=5.3U
M$19 vdd iref \$31 vdd pfet_03v3 L=2U W=2U AS=1.3P AD=0.52P PS=5.3U PD=2.52U
M$20 \$31 iref vdd vdd pfet_03v3 L=2U W=2U AS=0.52P AD=1.3P PS=2.52U PD=5.3U
M$21 GND \$4 \$4 GND nfet_03v3 L=2U W=2U AS=1.22P AD=0.52P PS=5.22U PD=2.52U
M$22 \$4 \$4 GND GND nfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$23 GND \$4 \$4 GND nfet_03v3 L=2U W=2U AS=0.52P AD=1.22P PS=2.52U PD=5.22U
M$24 \$5 \$4 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=0.52P PS=5.22U PD=2.52U
M$25 GND \$4 \$5 GND nfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$26 \$5 \$4 GND GND nfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$27 GND \$4 \$5 GND nfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$28 \$5 \$4 GND GND nfet_03v3 L=2U W=2U AS=0.52P AD=1.22P PS=2.52U PD=5.22U
M$29 GND \$5 \$5 GND nfet_03v3 L=1U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$30 PowerGate \$5 GND GND nfet_03v3 L=1U W=2U AS=1.22P AD=0.52P PS=5.22U
+ PD=2.52U
M$31 GND \$5 PowerGate GND nfet_03v3 L=1U W=2U AS=0.52P AD=0.52P PS=2.52U
+ PD=2.52U
M$32 PowerGate \$5 GND GND nfet_03v3 L=1U W=2U AS=0.52P AD=1.22P PS=2.52U
+ PD=5.22U
M$33 GND \$31 GND GND nfet_03v3 L=10U W=10U AS=6.1P AD=6.1P PS=21.22U PD=21.22U
M$34 GND \$31 GND GND nfet_03v3 L=10U W=10U AS=6.1P AD=6.1P PS=21.22U PD=21.22U
M$35 GND \$31 GND GND nfet_03v3 L=10U W=10U AS=6.1P AD=6.1P PS=21.22U PD=21.22U
M$36 GND \$31 GND GND nfet_03v3 L=10U W=10U AS=6.1P AD=6.1P PS=21.22U PD=21.22U
M$37 GND \$31 GND GND nfet_03v3 L=10U W=10U AS=6.1P AD=6.1P PS=21.22U PD=21.22U
M$38 GND \$31 GND GND nfet_03v3 L=10U W=10U AS=6.1P AD=6.1P PS=21.22U PD=21.22U
M$39 GND \$31 GND GND nfet_03v3 L=10U W=10U AS=6.1P AD=6.1P PS=21.22U PD=21.22U
M$40 GND \$31 GND GND nfet_03v3 L=10U W=10U AS=6.1P AD=6.1P PS=21.22U PD=21.22U
M$41 GND \$31 GND GND nfet_03v3 L=10U W=10U AS=6.1P AD=6.1P PS=21.22U PD=21.22U
.ENDS UndervoltageProtection
