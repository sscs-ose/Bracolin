* NGSPICE file created from PR_net.ext - technology: gf180mcuD

.subckt PR_net VSS VC VG_N IB_N VDD VB VA IB_P VG_P
X0 a_387_2075# VG_N.t0 VDD.t75 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1 VSS.t75 VSS.t74 VSS.t75 VSS.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2 VSS.t73 VSS.t72 VSS.t73 VSS.t9 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3 VDD.t71 VDD.t70 VDD.t71 VDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4 VSS.t71 VSS.t70 VSS.t71 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5 VSS.t69 VSS.t68 VSS.t69 VSS.t17 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6 VSS.t67 VSS.t66 VSS.t67 VSS.t3 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X7 VC VG_N.t1 a_387_151# VSS.t5 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X8 VDD.t69 VDD.t68 VDD.t69 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X9 a_375_8672# VG_P.t0 IB_P.t2 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X10 VSS.t65 VSS.t64 VSS.t65 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X11 VSS.t63 VSS.t62 VSS.t63 VSS.t9 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X12 VSS.t61 VSS.t60 VSS.t61 VSS.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X13 a_375_6740# VG_P.t1 VA.t0 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X14 VSS.t59 VSS.t58 VSS.t59 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X15 a_1781_8672# VG_P.t2 VSS.t1 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X16 a_1781_6740# VG_P.t3 a_n135_3233.t3 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X17 VSS.t57 VSS.t56 VSS.t57 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X18 VSS.t55 VSS.t54 VSS.t55 VSS.t3 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X19 VDD.t67 VDD.t66 VDD.t67 VDD.t25 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X20 VDD.t65 VDD.t64 VDD.t65 VDD.t25 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X21 VDD.t63 VDD.t61 VDD.t63 VDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X22 VSS.t53 VSS.t52 VSS.t53 VSS.t17 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X23 VSS.t51 VSS.t50 VSS.t51 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X24 VSS.t49 VSS.t48 VSS.t49 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X25 VDD.t60 VDD.t59 VDD.t60 VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X26 VSS.t47 VSS.t46 VSS.t47 VSS.t9 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X27 VSS.t45 VSS.t44 VSS.t45 VSS.t17 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X28 VDD.t58 VDD.t57 VDD.t58 VDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X29 VDD.t56 VDD.t55 VDD.t56 VDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X30 VDD.t54 VDD.t53 VDD.t54 VDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X31 VDD.t52 VDD.t51 VDD.t52 VDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X32 VDD VG_N.t2 a_1791_1309# VSS.t6 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X33 VDD.t50 VDD.t49 VDD.t50 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X34 VSS.t43 VSS.t42 VSS.t43 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X35 a_387_151# VG_N.t3 a_n135_151.t1 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X36 VSS.t41 VSS.t40 VSS.t41 VSS.t9 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X37 VSS.t39 VSS.t38 VSS.t39 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X38 VDD.t48 VDD.t47 VDD.t48 VDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X39 a_1791_151# VG_N.t4 VC.t0 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X40 VSS VG_P.t5 a_375_7906# VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X41 VA VG_P.t6 a_1781_9838# VDD.t6 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X42 VDD.t46 VDD.t45 VDD.t46 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X43 IB_P VG_P.t7 a_1781_7906# VDD.t6 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X44 VDD.t44 VDD.t43 VDD.t44 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X45 IB_N VG_N.t5 a_387_1309# VSS.t5 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X46 a_1791_1309# VG_N.t6 IB_N.t0 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X47 VDD.t42 VDD.t41 VDD.t42 VDD.t25 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X48 VDD.t40 VDD.t39 VDD.t40 VDD.t25 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X49 VSS.t37 VSS.t36 VSS.t37 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X50 a_387_1309# VG_N.t8 VDD.t74 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X51 VDD.t38 VDD.t37 VDD.t38 VDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X52 VDD.t36 VDD.t35 VDD.t36 VDD.t25 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X53 VSS.t35 VSS.t34 VSS.t35 VSS.t17 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X54 VDD.t34 VDD.t33 VDD.t34 VDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X55 VDD.t32 VDD.t31 VDD.t32 VDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X56 VDD.t30 VDD.t29 VDD.t30 VDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X57 VDD.t28 VDD.t27 VDD.t28 VDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X58 VDD.t26 VDD.t24 VDD.t26 VDD.t25 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X59 VDD VG_N.t10 a_1791_2075# VSS.t6 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X60 a_375_9838# VG_P.t8 VB.t0 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X61 a_375_7906# VG_P.t9 IB_P.t1 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X62 VSS.t33 VSS.t32 VSS.t33 VSS.t9 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X63 VDD.t23 VDD.t21 VDD.t23 VDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X64 VDD.t20 VDD.t18 VDD.t20 VDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X65 VC VG_N.t11 a_387_3233# VSS.t5 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X66 VSS.t31 VSS.t30 VSS.t31 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X67 a_1781_9838# VG_P.t10 a_n135_151.t3 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X68 a_1781_7906# VG_P.t11 VSS.t7 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X69 VDD.t17 VDD.t16 VDD.t17 VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X70 VSS VG_P.t12 a_375_8672# VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X71 VSS.t29 VSS.t28 VSS.t29 VSS.t6 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X72 a_1791_3233# VG_N.t12 VC.t2 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X73 VSS.t27 VSS.t26 VSS.t27 VSS.t17 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X74 VDD.t15 VDD.t14 VDD.t15 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X75 IB_P VG_P.t14 a_1781_8672# VDD.t6 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X76 VDD.t13 VDD.t12 VDD.t13 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X77 VB VG_P.t15 a_1781_6740# VDD.t6 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X78 VDD.t11 VDD.t10 VDD.t11 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X79 VSS.t25 VSS.t24 VSS.t25 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X80 IB_N VG_N.t13 a_387_2075# VSS.t5 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X81 VSS.t23 VSS.t21 VSS.t23 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X82 VSS.t20 VSS.t19 VSS.t20 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X83 a_387_3233# VG_N.t14 a_n135_3233.t1 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X84 VDD.t9 VDD.t8 VDD.t9 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X85 VSS.t18 VSS.t16 VSS.t18 VSS.t17 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X86 a_1791_2075# VG_N.t15 IB_N.t1 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X87 VSS.t15 VSS.t14 VSS.t15 VSS.t6 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X88 VDD.t7 VDD.t5 VDD.t7 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X89 VDD.t4 VDD.t2 VDD.t4 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X90 VSS.t13 VSS.t11 VSS.t13 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X91 VSS.t10 VSS.t8 VSS.t10 VSS.t9 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
R0 VG_N.n2 VG_N.t8 8.14051
R1 VG_N.n8 VG_N.t14 8.14051
R2 VG_N.n33 VG_N.t0 8.14051
R3 VG_N.n1 VG_N.t3 8.14051
R4 VG_N.n37 VG_N.t2 8.11137
R5 VG_N.n22 VG_N.t7 8.11137
R6 VG_N.n46 VG_N.t9 8.11137
R7 VG_N.n19 VG_N.t10 8.11137
R8 VG_N.n3 VG_N.t5 8.06917
R9 VG_N.n39 VG_N.t6 8.06917
R10 VG_N.n50 VG_N.t4 8.06917
R11 VG_N.n52 VG_N.t1 8.06917
R12 VG_N.n26 VG_N.t12 8.06917
R13 VG_N.n15 VG_N.t15 8.06917
R14 VG_N.n12 VG_N.t13 8.06917
R15 VG_N.n9 VG_N.t11 8.06917
R16 VG_N.n15 VG_N.n14 4.61892
R17 VG_N.n27 VG_N.n26 4.61892
R18 VG_N.n51 VG_N.n50 4.61892
R19 VG_N.n40 VG_N.n39 4.61892
R20 VG_N.n7 VG_N.n6 4.5005
R21 VG_N.n17 VG_N.n16 4.5005
R22 VG_N.n18 VG_N.n11 4.5005
R23 VG_N.n25 VG_N.n10 4.5005
R24 VG_N.n24 VG_N.n23 4.5005
R25 VG_N.n30 VG_N.n29 4.5005
R26 VG_N.n54 VG_N.n0 4.5005
R27 VG_N.n49 VG_N.n36 4.5005
R28 VG_N.n48 VG_N.n47 4.5005
R29 VG_N.n41 VG_N.n38 4.5005
R30 VG_N.n43 VG_N.n42 4.5005
R31 VG_N.n59 VG_N.n58 4.5005
R32 VG_N.n53 VG_N.n52 2.27692
R33 VG_N.n13 VG_N.n12 2.27692
R34 VG_N.n28 VG_N.n9 2.27692
R35 VG_N.n4 VG_N.n3 2.27692
R36 VG_N.n19 VG_N.n18 1.98105
R37 VG_N.n23 VG_N.n22 1.98105
R38 VG_N.n47 VG_N.n46 1.98105
R39 VG_N.n42 VG_N.n37 1.98105
R40 VG_N.n34 VG_N.n33 1.90721
R41 VG_N.n8 VG_N.n5 1.90721
R42 VG_N.n55 VG_N.n1 1.90721
R43 VG_N.n57 VG_N.n2 1.90721
R44 VG_N.n56 VG_N.n55 1.67168
R45 VG_N.n35 VG_N.n5 1.67138
R46 VG_N.n35 VG_N.n34 1.5005
R47 VG_N.n57 VG_N.n56 1.5005
R48 VG_N.n14 VG_N.n13 0.834997
R49 VG_N.n28 VG_N.n27 0.834997
R50 VG_N.n53 VG_N.n51 0.834997
R51 VG_N.n40 VG_N.n4 0.834997
R52 VG_N.n32 VG_N.n31 0.5099
R53 VG_N.n21 VG_N.n20 0.5099
R54 VG_N.n45 VG_N.n44 0.5099
R55 VG_N.n61 VG_N.n60 0.5099
R56 VG_N.n56 VG_N.n35 0.414926
R57 VG_N.n13 VG_N.n6 0.234207
R58 VG_N.n29 VG_N.n28 0.234207
R59 VG_N.n54 VG_N.n53 0.234207
R60 VG_N.n58 VG_N.n4 0.234207
R61 VG_N.n22 VG_N.n21 0.222597
R62 VG_N.n20 VG_N.n19 0.222597
R63 VG_N.n44 VG_N.n37 0.216676
R64 VG_N.n46 VG_N.n45 0.216676
R65 VG_N.n61 VG_N.n1 0.203347
R66 VG_N.n60 VG_N.n2 0.203347
R67 VG_N.n32 VG_N.n7 0.200632
R68 VG_N.n31 VG_N.n30 0.200632
R69 VG_N.n18 VG_N.n17 0.157683
R70 VG_N.n17 VG_N.n14 0.157683
R71 VG_N.n23 VG_N.n10 0.157683
R72 VG_N.n27 VG_N.n10 0.157683
R73 VG_N.n47 VG_N.n36 0.157683
R74 VG_N.n51 VG_N.n36 0.157683
R75 VG_N.n42 VG_N.n41 0.157683
R76 VG_N.n41 VG_N.n40 0.157683
R77 VG_N.n31 VG_N.n8 0.15361
R78 VG_N.n33 VG_N.n32 0.15361
R79 VG_N.n61 VG_N.n0 0.150895
R80 VG_N.n60 VG_N.n59 0.150895
R81 VG_N.n16 VG_N.n11 0.147342
R82 VG_N.n25 VG_N.n24 0.147342
R83 VG_N.n49 VG_N.n48 0.147342
R84 VG_N.n43 VG_N.n38 0.147342
R85 VG_N.n52 VG_N.n0 0.118921
R86 VG_N.n12 VG_N.n7 0.118921
R87 VG_N.n30 VG_N.n9 0.118921
R88 VG_N.n59 VG_N.n3 0.118921
R89 VG_N.n48 VG_N.n45 0.110632
R90 VG_N.n44 VG_N.n43 0.110632
R91 VG_N.n20 VG_N.n11 0.104711
R92 VG_N.n24 VG_N.n21 0.104711
R93 VG_N.n34 VG_N.n6 0.0474014
R94 VG_N.n29 VG_N.n5 0.0474014
R95 VG_N.n55 VG_N.n54 0.0474014
R96 VG_N.n58 VG_N.n57 0.0474014
R97 VG_N.n16 VG_N.n15 0.0289211
R98 VG_N.n26 VG_N.n25 0.0289211
R99 VG_N.n50 VG_N.n49 0.0289211
R100 VG_N.n39 VG_N.n38 0.0289211
R101 VG_N VG_N.n61 0.0131
R102 VDD.n60 VDD.n4 235.025
R103 VDD.n76 VDD.n4 234.572
R104 VDD.n76 VDD.n5 228.672
R105 VDD.n60 VDD.n5 225.946
R106 VDD.t25 VDD.t6 142.93
R107 VDD.t19 VDD.t62 142.93
R108 VDD.n47 VDD.n5 123.54
R109 VDD.n74 VDD.n4 117.733
R110 VDD.t3 VDD.t25 96.8792
R111 VDD.t6 VDD.t1 96.8792
R112 VDD.t62 VDD.t0 96.8792
R113 VDD.t22 VDD.t19 96.8792
R114 VDD.n76 VDD.t3 81.1238
R115 VDD.n60 VDD.t22 81.1238
R116 VDD.t1 VDD.n75 70.2717
R117 VDD.t0 VDD.n6 64.1315
R118 VDD.n75 VDD.n6 8.52856
R119 VDD.n11 VDD.t35 8.10567
R120 VDD.n11 VDD.t49 8.10567
R121 VDD.n0 VDD.t66 8.10567
R122 VDD.n0 VDD.t45 8.10567
R123 VDD.n79 VDD.t41 8.10567
R124 VDD.n79 VDD.t12 8.10567
R125 VDD.n28 VDD.t64 8.10567
R126 VDD.n28 VDD.t43 8.10567
R127 VDD.n29 VDD.t39 8.10567
R128 VDD.n29 VDD.t10 8.10567
R129 VDD.n32 VDD.t24 8.10567
R130 VDD.n32 VDD.t2 8.10567
R131 VDD.n69 VDD.t70 8.10567
R132 VDD.n18 VDD.t68 8.10567
R133 VDD.n7 VDD.t16 8.10567
R134 VDD.n14 VDD.t14 8.10567
R135 VDD.n66 VDD.t47 8.10567
R136 VDD.n66 VDD.t37 8.10567
R137 VDD.n64 VDD.t57 8.10567
R138 VDD.n64 VDD.t55 8.10567
R139 VDD.n63 VDD.t33 8.10567
R140 VDD.n63 VDD.t31 8.10567
R141 VDD.n58 VDD.t53 8.10567
R142 VDD.n58 VDD.t51 8.10567
R143 VDD.n57 VDD.t29 8.10567
R144 VDD.n57 VDD.t27 8.10567
R145 VDD.n55 VDD.t21 8.10567
R146 VDD.n55 VDD.t18 8.10567
R147 VDD.n25 VDD.t61 8.10567
R148 VDD.n50 VDD.t8 8.10567
R149 VDD.n26 VDD.t59 8.10567
R150 VDD.n43 VDD.t5 8.10567
R151 VDD.n41 VDD.n40 5.96085
R152 VDD.n40 VDD.n39 5.3195
R153 VDD.n42 VDD.n41 4.57315
R154 VDD.n41 VDD.n35 4.56231
R155 VDD.n39 VDD.t75 3.8555
R156 VDD.n38 VDD.n36 3.85313
R157 VDD.n38 VDD.n37 3.68497
R158 VDD.n39 VDD.t74 3.68261
R159 VDD.n68 VDD.t71 3.20383
R160 VDD.n72 VDD.t69 3.20383
R161 VDD.n17 VDD.t17 3.20383
R162 VDD.n13 VDD.t15 3.20383
R163 VDD.n53 VDD.t63 3.20383
R164 VDD.n49 VDD.t9 3.20383
R165 VDD.n46 VDD.t60 3.20383
R166 VDD.n27 VDD.t7 3.20383
R167 VDD.n45 VDD.n44 1.73383
R168 VDD.n52 VDD.n51 1.73383
R169 VDD.n16 VDD.n15 1.73383
R170 VDD.n71 VDD.n70 1.73383
R171 VDD.n40 VDD.n38 1.51393
R172 VDD.t69 VDD.n71 1.4705
R173 VDD.n71 VDD.t71 1.4705
R174 VDD.n16 VDD.t15 1.4705
R175 VDD.t17 VDD.n16 1.4705
R176 VDD.n52 VDD.t9 1.4705
R177 VDD.t63 VDD.n52 1.4705
R178 VDD.n45 VDD.t7 1.4705
R179 VDD.t60 VDD.n45 1.4705
R180 VDD.n8 VDD.t50 1.00929
R181 VDD.n9 VDD.t46 1.00929
R182 VDD.n1 VDD.t13 1.00929
R183 VDD.n2 VDD.t44 1.00929
R184 VDD.n30 VDD.t11 1.00929
R185 VDD.n33 VDD.t4 1.00929
R186 VDD.n19 VDD.t38 1.00929
R187 VDD.n20 VDD.t56 1.00929
R188 VDD.n21 VDD.t32 1.00929
R189 VDD.n22 VDD.t52 1.00929
R190 VDD.n23 VDD.t28 1.00929
R191 VDD.n24 VDD.t20 1.00929
R192 VDD.n8 VDD.t36 1.00871
R193 VDD.n9 VDD.t67 1.00871
R194 VDD.n1 VDD.t42 1.00871
R195 VDD.n2 VDD.t65 1.00871
R196 VDD.n30 VDD.t40 1.00871
R197 VDD.n33 VDD.t26 1.00871
R198 VDD.n19 VDD.t48 1.00871
R199 VDD.n20 VDD.t58 1.00871
R200 VDD.n21 VDD.t34 1.00871
R201 VDD.n22 VDD.t54 1.00871
R202 VDD.n23 VDD.t30 1.00871
R203 VDD.n24 VDD.t23 1.00871
R204 VDD.n54 VDD.n24 0.468749
R205 VDD.n56 VDD.n23 0.468749
R206 VDD.n59 VDD.n22 0.468749
R207 VDD.n62 VDD.n21 0.468749
R208 VDD.n65 VDD.n20 0.468749
R209 VDD.n67 VDD.n19 0.468749
R210 VDD.n34 VDD.n33 0.468749
R211 VDD.n31 VDD.n30 0.468749
R212 VDD.n3 VDD.n2 0.468749
R213 VDD.n78 VDD.n1 0.468749
R214 VDD.n10 VDD.n9 0.468749
R215 VDD.n12 VDD.n8 0.468749
R216 VDD.n61 VDD.n60 0.10728
R217 VDD.n74 VDD.n73 0.10728
R218 VDD.n75 VDD.n74 0.10728
R219 VDD.n77 VDD.n76 0.10728
R220 VDD.n48 VDD.n47 0.1055
R221 VDD.n47 VDD.n6 0.1055
R222 VDD.n66 VDD.n65 0.0382419
R223 VDD.n56 VDD.n55 0.0382419
R224 VDD.n11 VDD.n10 0.0382419
R225 VDD.n32 VDD.n31 0.0382419
R226 VDD.n64 VDD.n63 0.0364748
R227 VDD.n58 VDD.n57 0.0364748
R228 VDD.n29 VDD.n28 0.0364748
R229 VDD.n14 VDD.n13 0.0346711
R230 VDD.n15 VDD.n14 0.0346711
R231 VDD.n15 VDD.n7 0.0346711
R232 VDD.n17 VDD.n7 0.0346711
R233 VDD.n72 VDD.n18 0.0346711
R234 VDD.n70 VDD.n18 0.0346711
R235 VDD.n70 VDD.n69 0.0346711
R236 VDD.n69 VDD.n68 0.0346711
R237 VDD.n54 VDD.n53 0.0308563
R238 VDD.n68 VDD.n67 0.0308128
R239 VDD.n13 VDD.n12 0.0308128
R240 VDD.n44 VDD.n43 0.0293162
R241 VDD.n44 VDD.n26 0.0293162
R242 VDD.n46 VDD.n26 0.0293162
R243 VDD.n50 VDD.n49 0.0293162
R244 VDD.n51 VDD.n50 0.0293162
R245 VDD.n51 VDD.n25 0.0293162
R246 VDD.n53 VDD.n25 0.0293162
R247 VDD.n62 VDD.n61 0.0270708
R248 VDD.n78 VDD.n77 0.0270708
R249 VDD.n35 VDD.n34 0.0243625
R250 VDD.n43 VDD.n42 0.0232283
R251 VDD.n61 VDD.n59 0.0222742
R252 VDD.n77 VDD.n3 0.0222742
R253 VDD VDD.n0 0.0198759
R254 VDD.n67 VDD.n66 0.0193079
R255 VDD.n65 VDD.n64 0.0193079
R256 VDD.n63 VDD.n62 0.0193079
R257 VDD.n59 VDD.n58 0.0193079
R258 VDD.n57 VDD.n56 0.0193079
R259 VDD.n55 VDD.n54 0.0193079
R260 VDD.n12 VDD.n11 0.0193079
R261 VDD.n10 VDD.n0 0.0193079
R262 VDD.n79 VDD.n78 0.0193079
R263 VDD.n28 VDD.n3 0.0193079
R264 VDD.n31 VDD.n29 0.0193079
R265 VDD.n34 VDD.n32 0.0193079
R266 VDD.n48 VDD.n46 0.0185609
R267 VDD.n73 VDD.n72 0.0175856
R268 VDD VDD.n79 0.0170989
R269 VDD.n73 VDD.n17 0.0159011
R270 VDD.n49 VDD.n48 0.00983484
R271 VDD.n35 VDD.n27 0.0069938
R272 VDD.n42 VDD.n27 0.00658794
R273 VSS.t12 VSS.t6 401.067
R274 VSS.t4 VSS.t9 401.067
R275 VSS.t17 VSS.t12 273.233
R276 VSS.t6 VSS.t3 273.233
R277 VSS.t5 VSS.t4 273.233
R278 VSS.t9 VSS.t22 273.233
R279 VSS.n15 VSS.n5 250.45
R280 VSS.n67 VSS.n5 248.333
R281 VSS.n15 VSS.t17 227.945
R282 VSS.t22 VSS.n67 227.945
R283 VSS.t3 VSS.n6 196.143
R284 VSS.n36 VSS.n7 191.317
R285 VSS.n68 VSS.t5 191.263
R286 VSS.n67 VSS.n7 139.233
R287 VSS.n15 VSS.n7 138.493
R288 VSS.n69 VSS.n5 134.853
R289 VSS.n68 VSS.n6 24.3962
R290 VSS.n21 VSS.t64 8.06917
R291 VSS.n21 VSS.t52 8.06917
R292 VSS.n19 VSS.t24 8.06917
R293 VSS.n19 VSS.t16 8.06917
R294 VSS.n18 VSS.t11 8.06917
R295 VSS.n18 VSS.t68 8.06917
R296 VSS.n0 VSS.t36 8.06917
R297 VSS.n0 VSS.t34 8.06917
R298 VSS.n79 VSS.t19 8.06917
R299 VSS.n79 VSS.t26 8.06917
R300 VSS.n77 VSS.t50 8.06917
R301 VSS.n77 VSS.t44 8.06917
R302 VSS.n8 VSS.t58 8.06917
R303 VSS.n39 VSS.t74 8.06917
R304 VSS.n25 VSS.t66 8.06917
R305 VSS.n24 VSS.t28 8.06917
R306 VSS.n45 VSS.t42 8.06917
R307 VSS.n45 VSS.t46 8.06917
R308 VSS.n48 VSS.t70 8.06917
R309 VSS.n48 VSS.t72 8.06917
R310 VSS.n49 VSS.t56 8.06917
R311 VSS.n49 VSS.t62 8.06917
R312 VSS.n64 VSS.t30 8.06917
R313 VSS.n64 VSS.t32 8.06917
R314 VSS.n63 VSS.t21 8.06917
R315 VSS.n63 VSS.t8 8.06917
R316 VSS.n61 VSS.t38 8.06917
R317 VSS.n61 VSS.t40 8.06917
R318 VSS.n55 VSS.t48 8.06917
R319 VSS.n56 VSS.t60 8.06917
R320 VSS.n72 VSS.t54 8.06917
R321 VSS.n3 VSS.t14 8.06917
R322 VSS.n31 VSS.n30 7.29138
R323 VSS.n31 VSS.n9 4.57315
R324 VSS.n32 VSS.n31 4.56231
R325 VSS.n26 VSS.t7 3.73318
R326 VSS.n29 VSS.n28 3.73318
R327 VSS.n26 VSS.t1 3.4916
R328 VSS.n29 VSS.n27 3.4916
R329 VSS.n42 VSS.t59 3.3605
R330 VSS.n38 VSS.t75 3.3605
R331 VSS.n35 VSS.t67 3.3605
R332 VSS.n23 VSS.t29 3.3605
R333 VSS.n59 VSS.t49 3.3605
R334 VSS.t61 VSS.n4 3.3605
R335 VSS.n71 VSS.t55 3.3605
R336 VSS.n75 VSS.t15 3.3605
R337 VSS.n74 VSS.n73 2.1005
R338 VSS.n58 VSS.n57 2.1005
R339 VSS.n34 VSS.n33 2.1005
R340 VSS.n41 VSS.n40 2.1005
R341 VSS.n41 VSS.t75 1.2605
R342 VSS.t59 VSS.n41 1.2605
R343 VSS.n34 VSS.t29 1.2605
R344 VSS.t67 VSS.n34 1.2605
R345 VSS.n58 VSS.t61 1.2605
R346 VSS.t49 VSS.n58 1.2605
R347 VSS.t15 VSS.n74 1.2605
R348 VSS.n74 VSS.t55 1.2605
R349 VSS.n10 VSS.t53 0.918039
R350 VSS.n11 VSS.t18 0.918039
R351 VSS.n12 VSS.t69 0.918039
R352 VSS.n13 VSS.t35 0.918039
R353 VSS.n1 VSS.t27 0.918039
R354 VSS.n2 VSS.t45 0.918039
R355 VSS.n43 VSS.t47 0.918039
R356 VSS.n46 VSS.t73 0.918039
R357 VSS.n50 VSS.t63 0.918039
R358 VSS.n52 VSS.t33 0.918039
R359 VSS.n53 VSS.t10 0.918039
R360 VSS.n54 VSS.t41 0.918039
R361 VSS.n10 VSS.t65 0.91749
R362 VSS.n11 VSS.t25 0.91749
R363 VSS.n12 VSS.t13 0.91749
R364 VSS.n13 VSS.t37 0.91749
R365 VSS.n1 VSS.t20 0.91749
R366 VSS.n2 VSS.t51 0.91749
R367 VSS.n43 VSS.t43 0.91749
R368 VSS.n46 VSS.t71 0.91749
R369 VSS.n50 VSS.t57 0.91749
R370 VSS.n52 VSS.t31 0.91749
R371 VSS.n53 VSS.t23 0.91749
R372 VSS.n54 VSS.t39 0.91749
R373 VSS.n60 VSS.n54 0.582999
R374 VSS.n62 VSS.n53 0.582999
R375 VSS.n65 VSS.n52 0.582999
R376 VSS.n51 VSS.n50 0.582999
R377 VSS.n47 VSS.n46 0.582999
R378 VSS.n44 VSS.n43 0.582999
R379 VSS.n76 VSS.n2 0.582999
R380 VSS.n78 VSS.n1 0.582999
R381 VSS.n14 VSS.n13 0.582999
R382 VSS.n17 VSS.n12 0.582999
R383 VSS.n20 VSS.n11 0.582999
R384 VSS.n22 VSS.n10 0.582999
R385 VSS.n30 VSS.n29 0.174974
R386 VSS.n30 VSS.n26 0.130788
R387 VSS.n67 VSS.n66 0.0886356
R388 VSS.n37 VSS.n36 0.0886356
R389 VSS.n36 VSS.n6 0.0886356
R390 VSS.n16 VSS.n15 0.0886356
R391 VSS.n70 VSS.n69 0.0871667
R392 VSS.n69 VSS.n68 0.0871667
R393 VSS.n47 VSS.n45 0.0390622
R394 VSS.n62 VSS.n61 0.0390622
R395 VSS.n21 VSS.n20 0.0385696
R396 VSS.n78 VSS.n77 0.0385696
R397 VSS.n49 VSS.n48 0.0371211
R398 VSS.n64 VSS.n63 0.0371211
R399 VSS.n19 VSS.n18 0.0366533
R400 VSS.n24 VSS.n23 0.0341
R401 VSS.n33 VSS.n24 0.0341
R402 VSS.n39 VSS.n38 0.0341
R403 VSS.n40 VSS.n39 0.0341
R404 VSS.n40 VSS.n8 0.0341
R405 VSS.n42 VSS.n8 0.0341
R406 VSS.n35 VSS.n9 0.03362
R407 VSS.n60 VSS.n59 0.0302339
R408 VSS.n66 VSS.n51 0.0301981
R409 VSS.n76 VSS.n75 0.0301505
R410 VSS.n44 VSS.n42 0.0300328
R411 VSS.n23 VSS.n22 0.0299989
R412 VSS.n17 VSS.n16 0.0298187
R413 VSS.n75 VSS.n3 0.0294988
R414 VSS.n73 VSS.n3 0.0294988
R415 VSS.n73 VSS.n72 0.0294988
R416 VSS.n72 VSS.n71 0.0294988
R417 VSS.n56 VSS.n4 0.0294988
R418 VSS.n57 VSS.n56 0.0294988
R419 VSS.n57 VSS.n55 0.0294988
R420 VSS.n59 VSS.n55 0.0294988
R421 VSS VSS.n0 0.023495
R422 VSS.n66 VSS.n65 0.0203634
R423 VSS.n16 VSS.n14 0.0201097
R424 VSS.n38 VSS.n37 0.01994
R425 VSS.n33 VSS.n32 0.0197
R426 VSS.n45 VSS.n44 0.0196517
R427 VSS.n48 VSS.n47 0.0196517
R428 VSS.n51 VSS.n49 0.0196517
R429 VSS.n65 VSS.n64 0.0196517
R430 VSS.n63 VSS.n62 0.0196517
R431 VSS.n61 VSS.n60 0.0196517
R432 VSS.n22 VSS.n21 0.019407
R433 VSS.n20 VSS.n19 0.019407
R434 VSS.n18 VSS.n17 0.019407
R435 VSS.n14 VSS.n0 0.019407
R436 VSS.n79 VSS.n78 0.019407
R437 VSS.n77 VSS.n76 0.019407
R438 VSS.n71 VSS.n70 0.0183136
R439 VSS.n37 VSS.n35 0.01514
R440 VSS.n32 VSS.n25 0.0149
R441 VSS VSS.n79 0.0136583
R442 VSS.n70 VSS.n4 0.0120995
R443 VSS.n25 VSS.n9 0.00098
R444 VC.n2 VC.n1 9.84127
R445 VC.n1 VC.t2 4.1605
R446 VC.n2 VC.t0 4.15932
R447 VC.n1 VC.n0 4.15747
R448 VC VC.n3 3.57366
R449 VC VC.n2 0.583126
R450 VG_P.n33 VG_P.t0 8.17385
R451 VG_P.n2 VG_P.t9 8.17299
R452 VG_P.n1 VG_P.t1 8.17134
R453 VG_P.n8 VG_P.t8 8.16754
R454 VG_P.n19 VG_P.t14 8.15339
R455 VG_P.n43 VG_P.t7 8.15277
R456 VG_P.n46 VG_P.t15 8.15161
R457 VG_P.n22 VG_P.t6 8.14892
R458 VG_P.n3 VG_P.t5 8.10567
R459 VG_P.n39 VG_P.t11 8.10567
R460 VG_P.n26 VG_P.t10 8.10567
R461 VG_P.n15 VG_P.t2 8.10567
R462 VG_P.n12 VG_P.t12 8.10567
R463 VG_P.n9 VG_P.t4 8.10567
R464 VG_P.n52 VG_P.t13 8.10567
R465 VG_P.n50 VG_P.t3 8.10567
R466 VG_P.n15 VG_P.n14 4.62603
R467 VG_P.n39 VG_P.n38 4.6244
R468 VG_P.n51 VG_P.n50 4.62126
R469 VG_P.n27 VG_P.n26 4.61407
R470 VG_P.n7 VG_P.n6 4.5005
R471 VG_P.n17 VG_P.n16 4.5005
R472 VG_P.n18 VG_P.n11 4.5005
R473 VG_P.n25 VG_P.n10 4.5005
R474 VG_P.n24 VG_P.n23 4.5005
R475 VG_P.n30 VG_P.n29 4.5005
R476 VG_P.n54 VG_P.n0 4.5005
R477 VG_P.n49 VG_P.n36 4.5005
R478 VG_P.n48 VG_P.n47 4.5005
R479 VG_P.n42 VG_P.n37 4.5005
R480 VG_P.n41 VG_P.n40 4.5005
R481 VG_P.n59 VG_P.n58 4.5005
R482 VG_P.n13 VG_P.n12 2.26271
R483 VG_P.n4 VG_P.n3 2.26206
R484 VG_P.n53 VG_P.n52 2.26082
R485 VG_P.n28 VG_P.n9 2.25797
R486 VG_P.n23 VG_P.n22 1.97162
R487 VG_P.n47 VG_P.n46 1.97099
R488 VG_P.n19 VG_P.n18 1.97058
R489 VG_P.n43 VG_P.n42 1.97031
R490 VG_P.n8 VG_P.n5 1.9364
R491 VG_P.n55 VG_P.n1 1.93496
R492 VG_P.n57 VG_P.n2 1.93434
R493 VG_P.n34 VG_P.n33 1.93401
R494 VG_P.n35 VG_P.n5 1.67564
R495 VG_P.n56 VG_P.n55 1.67199
R496 VG_P.n35 VG_P.n34 1.5005
R497 VG_P.n57 VG_P.n56 1.5005
R498 VG_P.n14 VG_P.n13 0.834997
R499 VG_P.n38 VG_P.n4 0.834981
R500 VG_P.n53 VG_P.n51 0.83495
R501 VG_P.n28 VG_P.n27 0.834879
R502 VG_P.n32 VG_P.n31 0.5171
R503 VG_P.n21 VG_P.n20 0.5171
R504 VG_P.n45 VG_P.n44 0.5117
R505 VG_P.n61 VG_P.n60 0.5117
R506 VG_P.n56 VG_P.n35 0.415534
R507 VG_P.n20 VG_P.n19 0.235431
R508 VG_P.n29 VG_P.n28 0.234321
R509 VG_P.n54 VG_P.n53 0.234252
R510 VG_P.n58 VG_P.n4 0.234222
R511 VG_P.n13 VG_P.n6 0.234207
R512 VG_P.n44 VG_P.n43 0.219569
R513 VG_P.n46 VG_P.n45 0.214076
R514 VG_P.n22 VG_P.n21 0.213292
R515 VG_P.n33 VG_P.n32 0.207822
R516 VG_P.n60 VG_P.n2 0.193486
R517 VG_P.n61 VG_P.n1 0.188685
R518 VG_P.n31 VG_P.n8 0.188385
R519 VG_P.n18 VG_P.n17 0.157683
R520 VG_P.n17 VG_P.n14 0.157683
R521 VG_P.n23 VG_P.n10 0.157683
R522 VG_P.n27 VG_P.n10 0.157683
R523 VG_P.n47 VG_P.n36 0.157683
R524 VG_P.n51 VG_P.n36 0.157683
R525 VG_P.n42 VG_P.n41 0.157683
R526 VG_P.n41 VG_P.n38 0.157683
R527 VG_P.n60 VG_P.n59 0.154786
R528 VG_P.n61 VG_P.n0 0.15088
R529 VG_P.n16 VG_P.n11 0.147342
R530 VG_P.n40 VG_P.n37 0.145435
R531 VG_P.n32 VG_P.n7 0.144974
R532 VG_P.n49 VG_P.n48 0.141766
R533 VG_P.n25 VG_P.n24 0.133357
R534 VG_P.n12 VG_P.n7 0.133132
R535 VG_P.n59 VG_P.n3 0.131409
R536 VG_P.n31 VG_P.n30 0.131214
R537 VG_P.n52 VG_P.n0 0.128095
R538 VG_P.n30 VG_P.n9 0.1205
R539 VG_P.n44 VG_P.n37 0.113877
R540 VG_P.n48 VG_P.n45 0.111006
R541 VG_P.n20 VG_P.n11 0.102342
R542 VG_P.n24 VG_P.n21 0.0926429
R543 VG_P.n34 VG_P.n6 0.0220493
R544 VG_P.n29 VG_P.n5 0.0220493
R545 VG_P.n55 VG_P.n54 0.0220493
R546 VG_P.n58 VG_P.n57 0.0220493
R547 VG_P.n16 VG_P.n15 0.0218158
R548 VG_P.n40 VG_P.n39 0.021539
R549 VG_P.n50 VG_P.n49 0.0210063
R550 VG_P.n26 VG_P.n25 0.0197857
R551 VG_P VG_P.n61 0.0113
R552 IB_P.n2 IB_P.n1 7.55998
R553 IB_P.n1 IB_P.t2 3.65383
R554 IB_P.n2 IB_P.n0 3.65146
R555 IB_P.n1 IB_P.t1 3.57094
R556 IB_P IB_P.n3 3.44068
R557 IB_P IB_P.n2 0.133132
R558 VA VA.n0 16.7521
R559 VA VA.t0 3.52475
R560 a_n135_3233.n0 a_n135_3233.t3 10.6239
R561 a_n135_3233.n0 a_n135_3233.t1 10.3566
R562 a_n135_3233.n0 a_n135_3233.n1 10.0407
R563 a_n135_3233.n2 a_n135_3233.n0 9.63183
R564 a_n135_151.n0 a_n135_151.t1 10.6581
R565 a_n135_151.n0 a_n135_151.t3 10.1798
R566 a_n135_151.n2 a_n135_151.n0 9.78059
R567 a_n135_151.n0 a_n135_151.n1 9.34796
R568 IB_N.n3 IB_N.t0 3.84484
R569 IB_N.n2 IB_N.n1 3.84484
R570 IB_N.n2 IB_N.n0 3.69326
R571 IB_N IB_N.t1 3.64116
R572 IB_N.n3 IB_N.n2 0.31987
R573 IB_N IB_N.n3 0.0526053
R574 VB VB.t0 17.297
R575 VB VB.n0 3.46199
C0 a_1791_2075# VDD 0.035282f
C1 IB_P a_1781_8672# 0.033453f
C2 VB VG_P 2.79614f
C3 VA VDD 1.07535f
C4 VC a_387_151# 0.0284f
C5 VG_N a_1791_151# 0.130866f
C6 IB_N a_387_1309# 0.029151f
C7 VDD a_375_6740# 0.021515f
C8 a_387_2075# VG_N 0.158107f
C9 IB_N VC 0.126419f
C10 VG_N a_387_3233# 0.136838f
C11 VDD a_387_1309# 0.042519f
C12 VC VDD 0.214491f
C13 IB_P VB 0.418592f
C14 VA a_375_6740# 0.02829f
C15 a_387_2075# IB_N 0.042325f
C16 a_375_7906# VG_P 0.157264f
C17 VG_P a_375_9838# 0.139172f
C18 VG_P a_1781_7906# 0.131658f
C19 a_387_2075# VDD 0.029136f
C20 VG_P a_1781_6740# 0.130094f
C21 VB a_1781_8672# 0.010024f
C22 VG_P VDD 10.2564f
C23 VG_N a_1791_1309# 0.132223f
C24 a_375_7906# IB_P 0.041194f
C25 IB_P a_1781_7906# 0.04756f
C26 a_375_8672# VA 0.01182f
C27 VA VG_P 3.94561f
C28 VC a_1791_151# 0.0284f
C29 IB_P VDD 0.982546f
C30 IB_N a_1791_1309# 0.037867f
C31 a_1781_9838# VDD 0.021314f
C32 VG_P a_375_6740# 0.137881f
C33 VDD a_1791_1309# 0.042519f
C34 VG_N a_1791_3233# 0.130866f
C35 VC a_387_3233# 0.0284f
C36 IB_P VA 0.16048f
C37 a_1781_9838# VA 0.02829f
C38 VB a_375_9838# 0.02829f
C39 a_375_8672# VG_P 0.15726f
C40 VB a_1781_6740# 0.02829f
C41 VG_N a_387_151# 0.135524f
C42 VB VDD 1.39371f
C43 a_375_8672# IB_P 0.029183f
C44 IB_N VG_N 0.887499f
C45 VA VB 0.209375f
C46 VG_N VDD 0.917647f
C47 IB_P VG_P 0.796774f
C48 a_1781_9838# VG_P 0.132974f
C49 VC a_1791_3233# 0.0284f
C50 VDD a_375_9838# 0.021314f
C51 a_1791_2075# VG_N 0.132223f
C52 IB_N VDD 1.28862f
C53 VDD a_1781_6740# 0.021515f
C54 VG_P a_1781_8672# 0.1317f
C55 VG_N a_387_1309# 0.158104f
C56 a_375_7906# VA 0.01182f
C57 VC VG_N 1.75221f
C58 a_1791_2075# IB_N 0.057866f
.ends

