* Extracted by KLayout with GF180MCU LVS runset on : 29/11/2023 22:06

.SUBCKT FC_nfets_x2 D2 D1 S1 S2 G1 G2 B
M$1 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$2 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$4 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$7 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$8 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$9 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$10 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$11 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$12 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$13 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$14 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$15 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$16 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$17 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$18 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$19 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$20 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$21 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$22 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$23 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$24 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$25 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$26 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$27 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$28 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$29 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$30 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$31 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$32 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$33 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$34 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$35 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$36 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$37 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$38 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$39 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$40 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$41 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$42 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$43 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$44 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$45 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$46 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$47 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$48 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$49 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$50 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$51 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$52 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$53 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$54 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$55 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$56 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$57 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$58 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$59 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$60 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$61 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$62 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$63 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$64 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$65 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$66 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$67 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$68 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$69 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$70 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$71 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$72 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$73 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$74 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$75 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$76 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$77 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$78 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$79 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$80 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$81 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$82 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$83 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$84 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$85 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$86 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$87 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$88 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$89 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$90 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$91 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$92 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$93 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$94 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$95 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$96 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$97 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$98 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$99 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$100 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$101 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$102 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$103 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$104 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$105 S2 G2 D2 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$106 D2 G2 S2 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$107 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$108 D1 G1 S1 B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$109 S1 G1 D1 B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$110 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$111 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$112 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$113 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$114 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$115 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$116 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$117 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$118 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$119 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$120 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$121 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$122 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$123 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$124 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$125 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$126 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$127 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$128 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$129 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$130 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$131 B B B B nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$132 B B B B nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
.ENDS FC_nfets_x2
