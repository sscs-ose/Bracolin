* NGSPICE file created from FC_top.ext - technology: gf180mcuD

.subckt FC_top VP VN VOUT IREF AVSS AVDD
X0 AVDD.t1280 AVDD.t1279 AVDD.t1280 AVDD.t177 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1 AVSS.t282 AVSS.t281 AVSS.t282 AVSS.t46 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2 AVDD a_5396_n6451.t106 a_5396_8177.t87 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3 AVDD IREF.t45 a_n13990_8177.t267 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4 AVDD.t1278 AVDD.t1277 AVDD.t1278 AVDD.t110 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5 AVDD.t1276 AVDD.t1275 AVDD.t1276 AVDD.t373 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X6 AVDD IREF.t46 a_n13990_8177.t266 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X7 AVDD IREF.t47 a_n13990_8177.t265 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X8 VOUT a_n11317_n20927.t1 a_5396_9163.t131 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X9 AVDD IREF.t48 a_n13990_8177.t264 AVDD.t152 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X10 AVDD.t1274 AVDD.t1273 AVDD.t1274 AVDD.t121 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X11 AVDD IREF.t49 a_n13990_8177.t263 AVDD.t152 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X12 AVDD.t1272 AVDD.t1271 AVDD.t1272 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X13 AVDD.t1270 AVDD.t1269 AVDD.t1270 AVDD.t121 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X14 AVDD.t1268 AVDD.t1267 AVDD.t1268 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X15 AVDD.t1266 AVDD.t1265 AVDD.t1266 AVDD.t110 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X16 AVSS.t280 AVSS.t279 AVSS.t280 AVSS.t77 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X17 AVDD a_5396_n6451.t108 a_5396_9163.t87 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X18 AVDD.t1264 AVDD.t1263 AVDD.t1264 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X19 AVDD.t1262 AVDD.t1261 AVDD.t1262 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X20 AVDD IREF.t42 IREF.t43 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X21 AVDD.t1260 AVDD.t1259 AVDD.t1260 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X22 AVDD a_5396_n6451.t111 a_5396_9163.t84 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X23 AVDD IREF.t53 a_n13990_8177.t260 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X24 VOUT a_n11317_n20927.t1 a_5396_9163.t130 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X25 AVDD.t1258 AVDD.t1257 AVDD.t1258 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X26 AVSS.t278 AVSS.t277 AVSS.t278 AVSS.t4 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X27 AVSS.t276 AVSS.t275 AVSS.t276 AVSS.t52 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X28 AVDD IREF.t55 a_n11737_n14973.t29 AVDD.t810 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X29 AVDD.t1256 AVDD.t1255 AVDD.t1256 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X30 AVDD.t1254 AVDD.t1253 AVDD.t1254 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X31 AVDD.t1252 AVDD.t1251 AVDD.t1252 AVDD.t875 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X32 AVSS a_n11737_n14973.t30 a_n13990_n5465.t139 AVSS.t85 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X33 AVDD.t1250 AVDD.t1249 AVDD.t1250 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X34 AVDD.t1248 AVDD.t1247 AVDD.t1248 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X35 AVSS.t274 AVSS.t273 AVSS.t274 AVSS.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X36 a_n1533_n15598# a_n11317_n20927.t4 a_n2101_n15598# AVDD.t394 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X37 AVDD a_5396_n6451.t114 a_5396_9163.t83 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X38 AVDD.t1246 AVDD.t1245 AVDD.t1246 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X39 VOUT a_n11317_n20927.t1 a_5396_9163.t129 AVDD.t177 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X40 AVDD.t1244 AVDD.t1243 AVDD.t1244 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X41 AVDD IREF.t57 a_n11737_n15980.t20 AVDD.t810 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X42 AVDD.t1242 AVDD.t1241 AVDD.t1242 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X43 AVDD IREF.t59 a_n13990_8177.t257 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X44 AVSS.t272 AVSS.t271 AVSS.t272 AVSS.t28 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X45 AVDD.t1240 AVDD.t1239 AVDD.t1240 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X46 VOUT a_n11317_n20927.t1 a_5396_9163.t128 AVDD.t177 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X47 AVDD.t1238 AVDD.t1237 AVDD.t1238 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X48 AVDD.t1236 AVDD.t1235 AVDD.t1236 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X49 AVDD a_5396_n6451.t115 a_5396_8177.t83 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X50 AVDD.t1234 AVDD.t1233 AVDD.t1234 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X51 AVDD.t1232 AVDD.t1231 AVDD.t1232 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X52 AVDD a_5396_n6451.t117 a_5396_9163.t82 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X53 AVDD.t1230 AVDD.t1229 AVDD.t1230 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X54 AVDD a_5396_n6451.t118 a_5396_9163.t81 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X55 AVDD.t1228 AVDD.t1227 AVDD.t1228 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X56 AVDD.t1226 AVDD.t1225 AVDD.t1226 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X57 AVDD IREF.t61 a_n13990_8177.t255 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X58 AVDD IREF.t62 a_n13990_8177.t254 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X59 AVDD.t1224 AVDD.t1223 AVDD.t1224 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X60 AVDD.t1222 AVDD.t1221 AVDD.t1222 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X61 AVSS.t270 AVSS.t269 AVSS.t270 AVSS.t43 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X62 AVDD.t1220 AVDD.t1219 AVDD.t1220 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X63 AVDD.t1218 AVDD.t1217 AVDD.t1218 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X64 a_n1533_n16323# a_n11317_n20927.t1 a_n2101_n16323# AVDD.t394 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X65 AVSS.t268 AVSS.t267 AVSS.t268 AVSS.t235 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X66 VOUT a_n11317_n20927.t1 a_5396_9163.t127 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X67 AVDD.t1216 AVDD.t1215 AVDD.t1216 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X68 AVDD.t1214 AVDD.t1213 AVDD.t1214 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X69 AVDD IREF.t65 a_n13990_8177.t251 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X70 AVDD.t1212 AVDD.t1211 AVDD.t1212 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X71 AVDD.t1210 AVDD.t1209 AVDD.t1210 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X72 AVDD.t1208 AVDD.t1207 AVDD.t1208 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X73 IREF IREF.t40 AVDD.t1726 AVDD.t480 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X74 AVDD.t1206 AVDD.t1205 AVDD.t1206 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X75 AVDD.t1204 AVDD.t1203 AVDD.t1204 AVDD.t810 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X76 AVDD.t1202 AVDD.t1201 AVDD.t1202 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X77 AVDD IREF.t68 a_n13990_8177.t250 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X78 AVDD IREF.t69 a_n11737_n15980.t19 AVDD.t638 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X79 AVDD IREF.t70 a_n13990_8177.t249 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X80 VOUT a_n11317_n20927.t1 a_5396_9163.t126 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X81 AVDD.t1200 AVDD.t1199 AVDD.t1200 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X82 AVDD IREF.t71 a_n13990_8177.t248 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X83 AVDD a_5396_n6451.t122 a_5396_8177.t81 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X84 AVDD IREF.t72 a_n13990_8177.t247 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X85 AVDD IREF.t74 a_n13990_8177.t245 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X86 a_n2101_n15598# a_n11317_n20927.t4 a_n2631_n16323# AVDD.t328 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X87 AVDD.t1198 AVDD.t1197 AVDD.t1198 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X88 AVDD.t1196 AVDD.t1195 AVDD.t1196 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X89 AVDD.t1194 AVDD.t1193 AVDD.t1194 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X90 AVDD.t1192 AVDD.t1191 AVDD.t1192 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X91 AVDD IREF.t75 a_n13990_8177.t244 AVDD.t152 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X92 AVDD.t1190 AVDD.t1189 AVDD.t1190 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X93 AVDD.t1188 AVDD.t1187 AVDD.t1188 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X94 AVDD.t1186 AVDD.t1185 AVDD.t1186 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X95 AVDD a_5396_n6451.t123 a_5396_8177.t80 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X96 AVDD.t1184 AVDD.t1183 AVDD.t1184 AVDD.t264 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X97 AVDD.t1182 AVDD.t1181 AVDD.t1182 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X98 AVDD IREF.t77 a_n11737_n15980.t18 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X99 VOUT a_n11317_n20927.t1 a_5396_9163.t125 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X100 AVDD.t1180 AVDD.t1179 AVDD.t1180 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X101 IREF IREF.t38 AVDD.t1725 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X102 AVDD.t1178 AVDD.t1177 AVDD.t1178 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X103 AVDD.t1176 AVDD.t1175 AVDD.t1176 AVDD.t155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X104 AVSS.t266 AVSS.t265 AVSS.t266 AVSS.t31 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X105 AVDD IREF.t81 a_n13990_8177.t240 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X106 AVDD a_5396_n6451.t124 a_5396_8177.t79 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X107 AVDD.t1174 AVDD.t1173 AVDD.t1174 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X108 AVDD a_5396_n6451.t126 a_5396_9163.t77 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X109 AVDD a_5396_n6451.t127 a_5396_8177.t77 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X110 AVDD.t1172 AVDD.t1171 AVDD.t1172 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X111 AVDD.t1170 AVDD.t1169 AVDD.t1170 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X112 VOUT a_n11317_n20927.t1 a_5396_9163.t124 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X113 AVDD IREF.t82 a_n11737_n14973.t27 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X114 AVSS.t264 AVSS.t263 AVSS.t264 AVSS.t25 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X115 AVSS.t262 AVSS.t261 AVSS.t262 AVSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X116 AVSS.t260 AVSS.t259 AVSS.t260 AVSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X117 AVDD.t1168 AVDD.t1167 AVDD.t1168 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X118 AVDD IREF.t83 a_n11737_n14973.t26 AVDD.t282 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X119 a_n2101_n16323# a_n11317_n20927.t1 a_n2631_n16323# AVDD.t328 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X120 VOUT a_n11317_n20927.t1 a_5396_9163.t123 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X121 AVDD a_5396_n6451.t128 a_5396_8177.t76 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X122 AVSS a_n11737_n14973.t38 a_n13990_n6451.t51 AVSS.t55 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X123 a_n6139_n21443# a_n11737_n15980.t27 a_n6661_n21443# AVSS.t178 nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X124 AVDD.t1166 AVDD.t1165 AVDD.t1166 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X125 AVDD.t1164 AVDD.t1163 AVDD.t1164 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X126 AVDD.t1162 AVDD.t1161 AVDD.t1162 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X127 AVDD IREF.t84 a_n13990_8177.t239 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X128 AVSS a_n11737_n14973.t39 a_n13990_n6451.t52 AVSS.t114 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X129 AVDD.t1160 AVDD.t1159 AVDD.t1160 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X130 VOUT a_n11317_n20927.t1 a_5396_9163.t122 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X131 AVDD.t1158 AVDD.t1157 AVDD.t1158 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X132 AVSS.t258 AVSS.t257 AVSS.t258 AVSS.t222 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X133 VOUT a_n11317_n20927.t1 a_5396_9163.t121 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X134 AVDD.t1156 AVDD.t1155 AVDD.t1156 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X135 AVDD.t1154 AVDD.t1153 AVDD.t1154 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X136 AVDD.t1152 AVDD.t1151 AVDD.t1152 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X137 AVDD.t1150 AVDD.t1149 AVDD.t1150 AVDD.t13 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X138 AVDD a_5396_n6451.t132 a_5396_8177.t74 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X139 AVDD.t1148 AVDD.t1147 AVDD.t1148 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X140 AVDD.t1146 AVDD.t1145 AVDD.t1146 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X141 AVDD.t1144 AVDD.t1143 AVDD.t1144 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X142 VOUT a_n11317_n20927.t1 a_5396_9163.t120 AVDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X143 a_n1533_n17634# a_n11317_n20927.t1 a_n2101_n17634# AVDD.t394 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X144 AVDD.t1142 AVDD.t1141 AVDD.t1142 AVDD.t180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X145 AVSS.t256 AVSS.t255 AVSS.t256 AVSS.t31 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X146 AVDD.t1140 AVDD.t1139 AVDD.t1140 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X147 AVDD.t1138 AVDD.t1137 AVDD.t1138 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X148 AVDD.t1136 AVDD.t1135 AVDD.t1136 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X149 AVSS.t254 AVSS.t253 AVSS.t254 AVSS.t4 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X150 AVSS a_n11737_n14973.t40 a_n13990_n6451.t53 AVSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X151 AVDD.t1134 AVDD.t1133 AVDD.t1134 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X152 AVDD.t1132 AVDD.t1131 AVDD.t1132 AVDD.t373 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X153 AVDD.t1130 AVDD.t1129 AVDD.t1130 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X154 AVDD IREF.t86 a_n13990_8177.t237 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X155 AVDD.t1128 AVDD.t1127 AVDD.t1128 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X156 AVDD.t1126 AVDD.t1125 AVDD.t1126 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X157 AVDD a_5396_n6451.t133 a_5396_9163.t74 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X158 AVDD IREF.t87 a_n13990_8177.t236 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X159 AVDD.t1124 AVDD.t1123 AVDD.t1124 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X160 AVDD.t1122 AVDD.t1121 AVDD.t1122 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X161 AVDD.t1120 AVDD.t1119 AVDD.t1120 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X162 AVDD.t1118 AVDD.t1117 AVDD.t1118 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X163 AVSS.t252 AVSS.t251 AVSS.t252 AVSS.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X164 AVDD.t1116 AVDD.t1115 AVDD.t1116 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X165 AVDD.t1114 AVDD.t1113 AVDD.t1114 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X166 AVDD IREF.t88 a_n13990_8177.t235 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X167 AVDD.t1112 AVDD.t1111 AVDD.t1112 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X168 AVDD IREF.t36 IREF.t37 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X169 AVDD IREF.t34 IREF.t35 AVDD.t638 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X170 AVSS.t250 AVSS.t249 AVSS.t250 AVSS.t77 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X171 AVDD.t1110 AVDD.t1109 AVDD.t1110 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X172 AVDD.t1108 AVDD.t1107 AVDD.t1108 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X173 AVDD.t1106 AVDD.t1105 AVDD.t1106 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X174 AVDD.t1104 AVDD.t1103 AVDD.t1104 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X175 AVDD.t1102 AVDD.t1101 AVDD.t1102 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X176 AVDD.t1100 AVDD.t1099 AVDD.t1100 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X177 AVDD.t1098 AVDD.t1097 AVDD.t1098 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X178 AVDD.t1096 AVDD.t1095 AVDD.t1096 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X179 AVDD.t1094 AVDD.t1093 AVDD.t1094 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X180 AVDD.t1092 AVDD.t1091 AVDD.t1092 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X181 AVDD IREF.t90 a_n13990_8177.t233 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X182 AVDD.t1090 AVDD.t1089 AVDD.t1090 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X183 AVDD.t1088 AVDD.t1087 AVDD.t1088 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X184 AVDD.t1086 AVDD.t1085 AVDD.t1086 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X185 VOUT a_n11317_n20927.t1 a_5396_9163.t119 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X186 AVDD IREF.t92 a_n13990_8177.t232 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X187 AVSS.t248 AVSS.t247 AVSS.t248 AVSS.t138 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X188 AVDD.t1084 AVDD.t1083 AVDD.t1084 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X189 AVSS.t246 AVSS.t245 AVSS.t246 AVSS.t49 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X190 AVDD IREF.t93 a_n13990_8177.t231 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X191 VOUT a_n11317_n20927.t1 a_5396_9163.t118 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X192 AVDD.t1082 AVDD.t1081 AVDD.t1082 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X193 AVDD.t1080 AVDD.t1079 AVDD.t1080 AVDD.t130 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X194 AVDD.t1078 AVDD.t1077 AVDD.t1078 AVDD.t192 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X195 AVDD.t1076 AVDD.t1075 AVDD.t1076 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X196 AVDD.t1074 AVDD.t1073 AVDD.t1074 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X197 AVDD.t1072 AVDD.t1071 AVDD.t1072 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X198 AVDD.t1070 AVDD.t1069 AVDD.t1070 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X199 AVDD.t1068 AVDD.t1067 AVDD.t1068 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X200 AVDD.t1066 AVDD.t1065 AVDD.t1066 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X201 AVDD a_5396_n6451.t135 a_5396_9163.t73 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X202 AVDD.t1064 AVDD.t1063 AVDD.t1064 AVDD.t195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X203 AVSS.t244 AVSS.t243 AVSS.t244 AVSS.t201 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X204 VOUT a_n11317_n20927.t1 a_5396_9163.t117 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X205 AVSS.t242 AVSS.t241 AVSS.t242 AVSS.t133 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X206 AVDD.t1062 AVDD.t1061 AVDD.t1062 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X207 AVDD.t1060 AVDD.t1059 AVDD.t1060 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X208 AVSS.t240 AVSS.t239 AVSS.t240 AVSS.t37 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X209 AVDD.t1058 AVDD.t1057 AVDD.t1058 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X210 a_n2101_n17634# a_n11317_n20927.t1 a_n2631_n17634# AVDD.t328 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X211 AVDD.t1056 AVDD.t1055 AVDD.t1056 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X212 AVDD a_5396_n6451.t137 a_5396_8177.t72 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X213 AVDD.t1054 AVDD.t1053 AVDD.t1054 AVDD.t152 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X214 AVDD IREF.t96 a_n13990_8177.t228 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X215 IREF IREF.t32 AVDD.t1720 AVDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X216 AVDD.t1052 AVDD.t1051 AVDD.t1052 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X217 AVDD.t1050 AVDD.t1049 AVDD.t1050 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X218 AVDD.t1048 AVDD.t1047 AVDD.t1048 AVDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X219 AVDD a_5396_n6451.t138 a_5396_9163.t71 AVDD.t155 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X220 AVDD.t1046 AVDD.t1045 AVDD.t1046 AVDD.t135 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X221 AVDD.t1044 AVDD.t1043 AVDD.t1044 AVDD.t638 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X222 AVSS.t238 AVSS.t237 AVSS.t238 AVSS.t46 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X223 AVDD.t1042 AVDD.t1041 AVDD.t1042 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X224 AVDD.t1040 AVDD.t1039 AVDD.t1040 AVDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X225 AVDD a_5396_n6451.t140 a_5396_8177.t71 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X226 AVDD.t1038 AVDD.t1037 AVDD.t1038 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X227 AVDD.t1036 AVDD.t1035 AVDD.t1036 AVDD.t135 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X228 AVDD.t1034 AVDD.t1033 AVDD.t1034 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X229 IREF IREF.t30 AVDD.t1719 AVDD.t480 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X230 AVDD a_5396_n6451.t141 a_5396_8177.t70 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X231 AVDD.t1032 AVDD.t1031 AVDD.t1032 AVDD.t135 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X232 AVDD a_5396_n6451.t142 a_5396_9163.t69 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X233 VOUT a_n11317_n20927.t1 a_5396_9163.t116 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X234 AVDD a_5396_n6451.t144 a_5396_8177.t68 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X235 AVSS.t236 AVSS.t234 AVSS.t236 AVSS.t235 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X236 AVDD.t1030 AVDD.t1029 AVDD.t1030 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X237 AVDD IREF.t99 a_n13990_8177.t227 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X238 AVDD.t1028 AVDD.t1027 AVDD.t1028 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X239 AVDD.t1026 AVDD.t1025 AVDD.t1026 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X240 AVDD IREF.t100 a_n13990_8177.t226 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X241 a_n6139_n20820# a_n11737_n15980.t36 a_n6661_n21443# AVSS.t178 nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X242 AVDD.t1024 AVDD.t1023 AVDD.t1024 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X243 VOUT a_n11737_n15980.t37 a_n13990_n5465.t36 AVSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X244 AVSS a_n11737_n14973.t42 a_n13990_n6451.t19 AVSS.t43 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X245 AVDD.t1022 AVDD.t1021 AVDD.t1022 AVDD.t121 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X246 AVDD IREF.t101 a_n11737_n14973.t24 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X247 AVDD.t1020 AVDD.t1019 AVDD.t1020 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X248 AVSS.t233 AVSS.t232 AVSS.t233 AVSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X249 AVDD.t1018 AVDD.t1017 AVDD.t1018 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X250 AVDD.t1016 AVDD.t1015 AVDD.t1016 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X251 AVDD.t1014 AVDD.t1013 AVDD.t1014 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X252 AVDD.t1012 AVDD.t1011 AVDD.t1012 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X253 AVDD.t1010 AVDD.t1009 AVDD.t1010 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X254 AVDD IREF.t102 a_n13990_8177.t225 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X255 AVDD a_5396_n6451.t147 a_5396_9163.t66 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X256 AVDD.t1008 AVDD.t1007 AVDD.t1008 AVDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X257 AVDD IREF.t28 IREF.t29 AVDD.t282 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X258 AVDD a_5396_n6451.t148 a_5396_8177.t67 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X259 AVDD IREF.t103 a_n13990_8177.t224 AVDD.t238 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X260 AVDD.t1006 AVDD.t1005 AVDD.t1006 AVDD.t195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X261 AVDD.t1004 AVDD.t1003 AVDD.t1004 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X262 AVDD IREF.t104 a_n11737_n15980.t17 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X263 AVSS a_n11737_n14973.t43 a_n13990_n6451.t20 AVSS.t85 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X264 a_n965_n16909# a_n11317_n20927.t1 a_n1533_n16909# AVDD.t264 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X265 AVDD.t1002 AVDD.t1001 AVDD.t1002 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X266 AVDD.t1000 AVDD.t999 AVDD.t1000 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X267 AVDD.t998 AVDD.t997 AVDD.t998 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X268 AVDD.t996 AVDD.t995 AVDD.t996 AVDD.t92 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X269 AVDD a_5396_n6451.t149 a_5396_9163.t65 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X270 AVDD.t994 AVDD.t993 AVDD.t994 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X271 AVSS.t231 AVSS.t230 AVSS.t231 AVSS.t28 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X272 AVDD a_5396_n6451.t150 a_5396_8177.t66 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X273 AVSS.t229 AVSS.t228 AVSS.t229 AVSS.t31 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X274 AVDD IREF.t105 a_n13990_8177.t223 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X275 AVDD.t992 AVDD.t991 AVDD.t992 AVDD.t2 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X276 AVDD.t990 AVDD.t989 AVDD.t990 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X277 AVDD.t988 AVDD.t987 AVDD.t988 AVDD.t195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X278 AVDD IREF.t106 a_n13990_8177.t222 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X279 AVDD.t986 AVDD.t985 AVDD.t986 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X280 AVSS a_n11737_n14973.t6 a_n11737_n14973.t7 AVSS.t138 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X281 AVSS.t227 AVSS.t226 AVSS.t227 AVSS.t175 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X282 AVDD.t984 AVDD.t983 AVDD.t984 AVDD.t180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X283 AVSS.t225 AVSS.t224 AVSS.t225 AVSS.t172 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X284 AVDD.t982 AVDD.t981 AVDD.t982 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X285 AVDD.t980 AVDD.t979 AVDD.t980 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X286 AVSS a_n11737_n14973.t44 a_n13990_n5465.t24 AVSS.t114 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X287 VOUT a_n11317_n20927.t1 a_5396_9163.t115 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X288 AVDD.t978 AVDD.t977 AVDD.t978 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X289 AVDD.t976 AVDD.t975 AVDD.t976 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X290 AVDD.t974 AVDD.t973 AVDD.t974 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X291 AVDD.t972 AVDD.t971 AVDD.t972 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X292 AVDD.t970 AVDD.t969 AVDD.t970 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X293 AVSS.t223 AVSS.t221 AVSS.t223 AVSS.t222 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X294 AVDD.t968 AVDD.t967 AVDD.t968 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X295 AVDD.t966 AVDD.t965 AVDD.t966 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X296 AVSS a_n11737_n14973.t45 a_n13990_n5465.t15 AVSS.t25 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X297 AVSS a_n11737_n14973.t46 a_n13990_n6451.t12 AVSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X298 AVSS a_n11737_n14973.t47 a_n13990_n5465.t16 AVSS.t19 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X299 AVDD.t964 AVDD.t963 AVDD.t964 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X300 AVDD.t962 AVDD.t961 AVDD.t962 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X301 AVSS a_n11737_n14973.t48 a_n11317_n20927.t1 AVSS.t133 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X302 AVDD.t960 AVDD.t959 AVDD.t960 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X303 AVDD.t958 AVDD.t957 AVDD.t958 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X304 AVDD.t956 AVDD.t955 AVDD.t956 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X305 AVSS.t220 AVSS.t219 AVSS.t220 AVSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X306 AVSS.t218 AVSS.t217 AVSS.t218 AVSS.t2 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X307 AVDD.t954 AVDD.t953 AVDD.t954 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X308 AVDD.t952 AVDD.t951 AVDD.t952 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X309 VOUT a_n11317_n20927.t1 a_5396_9163.t114 AVDD.t110 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X310 AVDD.t950 AVDD.t949 AVDD.t950 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X311 AVDD a_5396_n6451.t156 a_5396_9163.t64 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X312 AVDD.t948 AVDD.t947 AVDD.t948 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X313 AVDD IREF.t113 a_n13990_8177.t218 AVDD.t152 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X314 AVDD.t946 AVDD.t945 AVDD.t946 AVDD.t130 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X315 VOUT a_n11317_n20927.t1 a_5396_9163.t113 AVDD.t110 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X316 AVDD.t944 AVDD.t943 AVDD.t944 AVDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X317 AVDD.t942 AVDD.t941 AVDD.t942 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X318 AVDD a_5396_n6451.t158 a_5396_9163.t62 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X319 AVDD.t940 AVDD.t939 AVDD.t940 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X320 AVDD.t938 AVDD.t937 AVDD.t938 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X321 AVDD.t936 AVDD.t935 AVDD.t936 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X322 AVDD.t934 AVDD.t933 AVDD.t934 AVDD.t177 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X323 AVSS.t216 AVSS.t215 AVSS.t216 AVSS.t52 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X324 AVSS a_n11737_n14973.t49 a_n13990_n5465.t7 AVSS.t43 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X325 AVDD.t932 AVDD.t931 AVDD.t932 AVDD.t13 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X326 AVDD IREF.t116 a_n13990_8177.t215 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X327 AVDD.t930 AVDD.t929 AVDD.t930 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X328 AVDD IREF.t117 a_n13990_8177.t214 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X329 AVSS.t214 AVSS.t213 AVSS.t214 AVSS.t82 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X330 AVSS.t212 AVSS.t211 AVSS.t212 AVSS.t34 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X331 AVDD IREF.t119 a_n13990_8177.t212 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X332 AVSS.t210 AVSS.t209 AVSS.t210 AVSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X333 AVDD.t928 AVDD.t927 AVDD.t928 AVDD.t155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X334 AVDD.t926 AVDD.t925 AVDD.t926 AVDD.t27 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X335 AVDD.t924 AVDD.t923 AVDD.t924 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X336 AVDD.t922 AVDD.t921 AVDD.t922 AVDD.t92 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X337 AVDD a_5396_n6451.t160 a_5396_8177.t59 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X338 AVDD.t920 AVDD.t919 AVDD.t920 AVDD.t373 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X339 AVSS.t208 AVSS.t207 AVSS.t208 AVSS.t158 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X340 AVSS.t206 AVSS.t205 AVSS.t206 AVSS.t155 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X341 AVSS.t204 AVSS.t203 AVSS.t204 AVSS.t49 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X342 AVDD.t918 AVDD.t917 AVDD.t918 AVDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X343 AVDD.t916 AVDD.t915 AVDD.t916 AVDD.t110 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X344 AVDD.t914 AVDD.t913 AVDD.t914 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X345 AVDD.t912 AVDD.t911 AVDD.t912 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X346 AVDD.t910 AVDD.t909 AVDD.t910 AVDD.t92 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X347 AVDD.t908 AVDD.t907 AVDD.t908 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X348 AVDD.t906 AVDD.t905 AVDD.t906 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X349 AVDD.t904 AVDD.t903 AVDD.t904 AVDD.t92 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X350 AVSS.t202 AVSS.t200 AVSS.t202 AVSS.t201 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X351 AVSS.t199 AVSS.t198 AVSS.t199 AVSS.t70 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X352 AVSS.t197 AVSS.t196 AVSS.t197 AVSS.t67 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X353 AVDD.t902 AVDD.t901 AVDD.t902 AVDD.t480 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X354 IREF IREF.t26 AVDD.t1716 AVDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X355 AVDD.t900 AVDD.t899 AVDD.t900 AVDD.t92 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X356 AVSS a_n11737_n14973.t50 a_n13990_n5465.t8 AVSS.t55 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X357 AVDD.t898 AVDD.t897 AVDD.t898 AVDD.t13 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X358 VOUT a_n11317_n20927.t1 a_5396_9163.t112 AVDD.t192 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X359 AVDD a_5396_n6451.t164 a_5396_8177.t57 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X360 AVDD.t896 AVDD.t895 AVDD.t896 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X361 AVSS.t195 AVSS.t194 AVSS.t195 AVSS.t46 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X362 AVDD.t894 AVDD.t893 AVDD.t894 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X363 AVDD.t892 AVDD.t891 AVDD.t892 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X364 AVDD a_5396_n6451.t165 a_5396_9163.t59 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X365 AVDD.t890 AVDD.t889 AVDD.t890 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X366 AVDD a_5396_n6451.t166 a_5396_9163.t58 AVDD.t155 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X367 AVDD a_5396_n6451.t167 a_5396_8177.t56 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X368 AVDD IREF.t123 a_n11737_n14973.t21 AVDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X369 AVDD.t888 AVDD.t887 AVDD.t888 AVDD.t373 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X370 VOUT a_n11317_n20927.t1 a_5396_9163.t111 AVDD.t192 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X371 AVDD.t886 AVDD.t885 AVDD.t886 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X372 AVDD IREF.t124 a_n13990_8177.t209 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X373 AVDD.t884 AVDD.t883 AVDD.t884 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X374 AVSS.t193 AVSS.t192 AVSS.t193 AVSS.t37 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X375 AVDD.t882 AVDD.t881 AVDD.t882 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X376 AVDD.t880 AVDD.t879 AVDD.t880 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X377 AVDD.t878 AVDD.t877 AVDD.t878 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X378 AVSS a_n11737_n14973.t53 a_n13990_n5465.t21 AVSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X379 VOUT a_n11737_n15980.t41 a_n13990_n5465.t35 AVSS.t16 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X380 VOUT a_n11737_n15980.t42 a_n13990_n5465.t34 AVSS.t13 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X381 AVDD.t876 AVDD.t874 AVDD.t876 AVDD.t875 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X382 AVDD.t873 AVDD.t872 AVDD.t873 AVDD.t177 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X383 AVSS.t191 AVSS.t190 AVSS.t191 AVSS.t144 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X384 AVSS.t189 AVSS.t188 AVSS.t189 AVSS.t141 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X385 AVDD.t871 AVDD.t870 AVDD.t871 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X386 AVDD.t869 AVDD.t868 AVDD.t869 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X387 AVDD IREF.t126 a_n11737_n14973.t20 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X388 AVDD.t867 AVDD.t866 AVDD.t867 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X389 AVDD.t865 AVDD.t864 AVDD.t865 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X390 AVDD.t863 AVDD.t862 AVDD.t863 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X391 AVDD.t861 AVDD.t860 AVDD.t861 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X392 AVDD a_5396_n6451.t170 a_5396_8177.t54 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X393 AVSS.t187 AVSS.t186 AVSS.t187 AVSS.t178 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X394 AVDD.t859 AVDD.t858 AVDD.t859 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X395 AVDD.t857 AVDD.t856 AVDD.t857 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X396 AVDD.t855 AVDD.t854 AVDD.t855 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X397 AVDD IREF.t24 IREF.t25 AVDD.t282 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X398 AVDD.t853 AVDD.t852 AVDD.t853 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X399 AVDD.t851 AVDD.t850 AVDD.t851 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X400 AVDD.t849 AVDD.t848 AVDD.t849 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X401 AVSS a_n11737_n14973.t55 a_n13990_n5465.t22 AVSS.t85 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X402 AVDD.t847 AVDD.t846 AVDD.t847 AVDD.t192 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X403 AVDD.t845 AVDD.t844 AVDD.t845 AVDD.t177 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X404 AVDD.t843 AVDD.t842 AVDD.t843 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X405 AVDD.t841 AVDD.t840 AVDD.t841 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X406 AVDD.t839 AVDD.t838 AVDD.t839 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X407 AVDD a_5396_n6451.t173 a_5396_8177.t53 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X408 AVDD.t837 AVDD.t836 AVDD.t837 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X409 AVDD.t835 AVDD.t834 AVDD.t835 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X410 AVDD.t833 AVDD.t832 AVDD.t833 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X411 AVDD.t831 AVDD.t830 AVDD.t831 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X412 AVDD.t829 AVDD.t828 AVDD.t829 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X413 AVDD.t827 AVDD.t826 AVDD.t827 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X414 AVSS.t185 AVSS.t184 AVSS.t185 AVSS.t28 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X415 AVDD.t825 AVDD.t824 AVDD.t825 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X416 AVDD.t823 AVDD.t822 AVDD.t823 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X417 AVDD IREF.t134 a_n13990_8177.t200 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X418 AVDD.t821 AVDD.t820 AVDD.t821 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X419 AVDD a_5396_n6451.t174 a_5396_9163.t54 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X420 AVDD.t819 AVDD.t818 AVDD.t819 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X421 AVDD.t817 AVDD.t816 AVDD.t817 AVDD.t180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X422 AVSS.t183 AVSS.t182 AVSS.t183 AVSS.t82 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X423 AVDD.t815 AVDD.t814 AVDD.t815 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X424 IREF IREF.t22 AVDD.t1713 AVDD.t39 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X425 AVDD IREF.t138 a_n13990_8177.t198 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X426 AVDD a_5396_n6451.t176 a_5396_9163.t53 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X427 AVSS.t181 AVSS.t180 AVSS.t181 AVSS.t96 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X428 AVDD.t813 AVDD.t812 AVDD.t813 AVDD.t152 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X429 AVDD.t811 AVDD.t809 AVDD.t811 AVDD.t810 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X430 AVDD.t808 AVDD.t807 AVDD.t808 AVDD.t2 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X431 AVSS.t179 AVSS.t177 AVSS.t179 AVSS.t178 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X432 AVDD.t806 AVDD.t805 AVDD.t806 AVDD.t13 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X433 AVSS.t176 AVSS.t174 AVSS.t176 AVSS.t175 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X434 AVSS.t173 AVSS.t171 AVSS.t173 AVSS.t172 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X435 VOUT a_n11317_n20927.t1 a_5396_9163.t110 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X436 AVDD.t804 AVDD.t803 AVDD.t804 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X437 a_n965_n15598# a_n11317_n20927.t1 a_n1533_n15598# AVDD.t264 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X438 AVDD.t802 AVDD.t801 AVDD.t802 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X439 AVDD.t800 AVDD.t799 AVDD.t800 AVDD.t135 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X440 AVDD.t798 AVDD.t797 AVDD.t798 AVDD.t373 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X441 AVDD.t796 AVDD.t795 AVDD.t796 AVDD.t155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X442 AVDD.t794 AVDD.t793 AVDD.t794 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X443 AVDD IREF.t143 a_n13990_8177.t195 AVDD.t152 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X444 AVDD a_5396_n6451.t179 a_5396_9163.t52 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X445 AVDD.t792 AVDD.t791 AVDD.t792 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X446 AVDD.t790 AVDD.t789 AVDD.t790 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X447 AVDD.t788 AVDD.t787 AVDD.t788 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X448 AVDD IREF.t144 a_n13990_8177.t194 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X449 AVDD.t786 AVDD.t785 AVDD.t786 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X450 VOUT a_n11317_n20927.t1 a_5396_9163.t109 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X451 AVSS.t170 AVSS.t169 AVSS.t170 AVSS.t77 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X452 AVDD.t784 AVDD.t783 AVDD.t784 AVDD.t130 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X453 AVDD.t782 AVDD.t781 AVDD.t782 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X454 AVDD a_5396_n6451.t182 a_5396_9163.t50 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X455 AVDD.t780 AVDD.t779 AVDD.t780 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X456 AVDD.t778 AVDD.t777 AVDD.t778 AVDD.t121 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X457 AVDD.t776 AVDD.t775 AVDD.t776 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X458 VOUT a_n11317_n20927.t1 a_5396_9163.t108 AVDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X459 AVDD.t774 AVDD.t773 AVDD.t774 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X460 AVDD.t772 AVDD.t771 AVDD.t772 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X461 AVDD IREF.t147 a_n11737_n15980.t13 AVDD.t810 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X462 AVDD IREF.t149 a_n13990_8177.t190 AVDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X463 AVDD IREF.t150 a_n13990_8177.t189 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X464 AVDD.t770 AVDD.t769 AVDD.t770 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X465 AVDD.t768 AVDD.t767 AVDD.t768 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X466 AVDD.t766 AVDD.t765 AVDD.t766 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X467 AVDD.t764 AVDD.t763 AVDD.t764 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X468 a_n965_n16909# a_n11317_n20927.t1 a_n1533_n16323# AVDD.t264 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X469 AVSS.t168 AVSS.t167 AVSS.t168 AVSS.t52 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X470 AVDD.t762 AVDD.t761 AVDD.t762 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X471 AVDD IREF.t151 a_n11737_n14973.t18 AVDD.t282 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X472 AVDD IREF.t152 a_n13990_8177.t188 AVDD.t152 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X473 AVDD.t760 AVDD.t759 AVDD.t760 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X474 AVDD.t758 AVDD.t757 AVDD.t758 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X475 AVDD.t756 AVDD.t755 AVDD.t756 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X476 AVDD.t754 AVDD.t753 AVDD.t754 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X477 AVDD.t752 AVDD.t751 AVDD.t752 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X478 AVDD.t750 AVDD.t749 AVDD.t750 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X479 AVSS a_n11737_n14973.t58 a_n13990_n5465.t27 AVSS.t235 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X480 AVSS.t166 AVSS.t165 AVSS.t166 AVSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X481 AVSS.t164 AVSS.t162 AVSS.t164 AVSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X482 AVDD.t748 AVDD.t747 AVDD.t748 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X483 AVDD.t746 AVDD.t745 AVDD.t746 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X484 AVDD.t744 AVDD.t743 AVDD.t744 AVDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X485 AVDD a_5396_n6451.t185 a_5396_9163.t49 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X486 AVDD.t742 AVDD.t741 AVDD.t742 AVDD.t394 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X487 AVDD.t740 AVDD.t739 AVDD.t740 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X488 AVDD.t738 AVDD.t737 AVDD.t738 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X489 AVSS.t161 AVSS.t160 AVSS.t161 AVSS.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X490 AVSS.t159 AVSS.t157 AVSS.t159 AVSS.t158 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X491 AVDD.t736 AVDD.t735 AVDD.t736 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X492 AVDD.t734 AVDD.t733 AVDD.t734 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X493 AVSS.t156 AVSS.t154 AVSS.t156 AVSS.t155 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X494 AVDD IREF.t155 a_n11737_n15980.t12 AVDD.t282 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X495 AVSS.t153 AVSS.t152 AVSS.t153 AVSS.t16 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X496 AVSS.t151 AVSS.t150 AVSS.t151 AVSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X497 AVSS.t149 AVSS.t148 AVSS.t149 AVSS.t37 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X498 AVDD.t732 AVDD.t731 AVDD.t732 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X499 AVSS a_n11737_n15980.t44 a_n6139_n21443# AVSS.t99 nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X500 AVDD.t730 AVDD.t729 AVDD.t730 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X501 AVDD.t728 AVDD.t727 AVDD.t728 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X502 AVSS a_n11737_n14973.t60 a_n13990_n6451.t24 AVSS.t55 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X503 AVDD.t726 AVDD.t725 AVDD.t726 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X504 AVDD.t724 AVDD.t723 AVDD.t724 AVDD.t180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X505 AVDD.t722 AVDD.t721 AVDD.t722 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X506 AVDD.t720 AVDD.t719 AVDD.t720 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X507 AVDD.t718 AVDD.t716 AVDD.t718 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X508 AVDD.t715 AVDD.t714 AVDD.t715 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X509 AVDD.t713 AVDD.t712 AVDD.t713 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X510 AVDD.t711 AVDD.t710 AVDD.t711 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X511 AVDD.t709 AVDD.t708 AVDD.t709 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X512 AVDD.t707 AVDD.t706 AVDD.t707 AVDD.t180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X513 AVDD.t705 AVDD.t704 AVDD.t705 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X514 AVDD IREF.t20 IREF.t21 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X515 AVDD IREF.t159 a_n13990_8177.t182 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X516 AVDD.t703 AVDD.t702 AVDD.t703 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X517 AVDD.t701 AVDD.t700 AVDD.t701 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X518 AVDD.t699 AVDD.t698 AVDD.t699 AVDD.t192 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X519 AVDD IREF.t160 a_n13990_8177.t181 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X520 AVDD.t697 AVDD.t696 AVDD.t697 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X521 AVDD.t695 AVDD.t694 AVDD.t695 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X522 AVDD.t693 AVDD.t692 AVDD.t693 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X523 AVDD.t691 AVDD.t690 AVDD.t691 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X524 AVDD.t689 AVDD.t688 AVDD.t689 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X525 AVDD.t687 AVDD.t686 AVDD.t687 AVDD.t282 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X526 AVDD.t685 AVDD.t684 AVDD.t685 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X527 AVDD.t683 AVDD.t682 AVDD.t683 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X528 AVDD a_5396_n6451.t190 a_5396_8177.t44 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X529 VOUT a_n11317_n20927.t1 a_5396_9163.t107 AVDD.t155 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X530 AVDD a_5396_n6451.t191 a_5396_9163.t46 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X531 AVSS.t147 AVSS.t146 AVSS.t147 AVSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X532 AVDD.t681 AVDD.t680 AVDD.t681 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X533 AVDD.t679 AVDD.t678 AVDD.t679 AVDD.t130 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X534 AVDD.t677 AVDD.t676 AVDD.t677 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X535 AVSS.t145 AVSS.t143 AVSS.t145 AVSS.t144 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X536 AVSS.t142 AVSS.t140 AVSS.t142 AVSS.t141 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X537 AVDD.t675 AVDD.t674 AVDD.t675 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X538 AVDD.t673 AVDD.t672 AVDD.t673 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X539 AVDD.t671 AVDD.t670 AVDD.t671 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X540 AVDD.t669 AVDD.t668 AVDD.t669 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X541 AVDD.t667 AVDD.t666 AVDD.t667 AVDD.t328 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X542 AVDD IREF.t162 a_n13990_8177.t179 AVDD.t152 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X543 AVDD a_5396_n6451.t193 a_5396_9163.t45 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X544 AVDD IREF.t163 a_n13990_8177.t178 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X545 AVDD a_5396_n6451.t194 a_5396_8177.t42 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X546 AVDD.t665 AVDD.t664 AVDD.t665 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X547 AVDD IREF.t164 a_n13990_8177.t177 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X548 AVDD.t663 AVDD.t662 AVDD.t663 AVDD.t152 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X549 AVDD a_5396_n6451.t195 a_5396_8177.t41 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X550 AVSS a_n11737_n14973.t63 a_n13990_n6451.t10 AVSS.t43 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X551 AVDD.t661 AVDD.t660 AVDD.t661 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X552 AVSS a_n11737_n14973.t64 a_n13990_n6451.t11 AVSS.t222 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X553 AVDD.t659 AVDD.t658 AVDD.t659 AVDD.t130 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X554 AVDD a_5396_n6451.t197 a_5396_9163.t43 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X555 AVDD a_n11317_n20927.t1 a_n1533_n17634# AVDD.t264 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X556 AVDD.t657 AVDD.t656 AVDD.t657 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X557 AVDD.t655 AVDD.t654 AVDD.t655 AVDD.t180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X558 VOUT a_n11317_n20927.t1 a_5396_9163.t106 AVDD.t177 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X559 AVDD.t653 AVDD.t652 AVDD.t653 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X560 AVDD.t651 AVDD.t650 AVDD.t651 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X561 AVSS.t139 AVSS.t137 AVSS.t139 AVSS.t138 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X562 a_n6139_n20267# a_n11737_n15980.t0 a_n11737_n15980.t1 AVSS.t178 nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X563 AVDD.t649 AVDD.t648 AVDD.t649 AVDD.t110 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X564 AVDD.t647 AVDD.t646 AVDD.t647 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X565 AVDD.t645 AVDD.t644 AVDD.t645 AVDD.t135 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X566 AVDD.t643 AVDD.t642 AVDD.t643 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X567 AVDD.t641 AVDD.t640 AVDD.t641 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X568 AVDD.t639 AVDD.t637 AVDD.t639 AVDD.t638 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X569 AVDD.t636 AVDD.t635 AVDD.t636 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X570 AVDD.t634 AVDD.t633 AVDD.t634 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X571 VOUT a_n11317_n20927.t1 a_5396_9163.t105 AVDD.t177 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X572 IREF IREF.t18 AVDD.t1710 AVDD.t39 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X573 AVSS.t136 AVSS.t135 AVSS.t136 AVSS.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X574 VOUT a_n11317_n20927.t1 a_5396_9163.t104 AVDD.t192 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X575 AVDD.t632 AVDD.t631 AVDD.t632 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X576 AVSS.t134 AVSS.t132 AVSS.t134 AVSS.t133 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X577 AVDD.t630 AVDD.t629 AVDD.t630 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X578 AVDD.t628 AVDD.t627 AVDD.t628 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X579 AVDD a_5396_n6451.t198 a_5396_9163.t42 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X580 AVSS.t131 AVSS.t130 AVSS.t131 AVSS.t114 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X581 AVDD.t626 AVDD.t625 AVDD.t626 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X582 AVDD.t624 AVDD.t623 AVDD.t624 AVDD.t121 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X583 AVDD.t622 AVDD.t621 AVDD.t622 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X584 AVDD.t620 AVDD.t619 AVDD.t620 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X585 VOUT a_n11317_n20927.t1 a_5396_9163.t103 AVDD.t192 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X586 AVDD a_5396_n6451.t201 a_5396_8177.t39 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X587 AVDD.t618 AVDD.t617 AVDD.t618 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X588 AVDD a_5396_n6451.t202 a_5396_9163.t40 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X589 VOUT a_n11317_n20927.t1 a_5396_9163.t102 AVDD.t155 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X590 AVDD IREF.t174 a_n13990_8177.t169 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X591 AVDD.t616 AVDD.t615 AVDD.t616 AVDD.t130 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X592 AVDD.t614 AVDD.t613 AVDD.t614 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X593 AVDD.t612 AVDD.t611 AVDD.t612 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X594 AVDD.t610 AVDD.t609 AVDD.t610 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X595 AVDD.t608 AVDD.t607 AVDD.t608 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X596 AVDD.t606 AVDD.t605 AVDD.t606 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X597 AVDD.t604 AVDD.t603 AVDD.t604 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X598 AVDD.t602 AVDD.t601 AVDD.t602 AVDD.t195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X599 AVDD.t600 AVDD.t599 AVDD.t600 AVDD.t152 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X600 AVDD.t598 AVDD.t597 AVDD.t598 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X601 AVSS a_n11737_n14973.t67 a_n13990_n6451.t3 AVSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X602 AVDD IREF.t175 a_n11737_n14973.t16 AVDD.t638 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X603 AVDD.t596 AVDD.t595 AVDD.t596 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X604 AVSS a_n11737_n14973.t68 a_n13990_n5465.t5 AVSS.t201 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X605 AVDD.t594 AVDD.t593 AVDD.t594 AVDD.t152 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X606 AVDD.t592 AVDD.t591 AVDD.t592 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X607 AVDD IREF.t177 a_n13990_8177.t167 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X608 a_n5579_n20820# a_n11737_n15980.t48 a_n6139_n20820# AVSS.t99 nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X609 AVDD.t590 AVDD.t589 AVDD.t590 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X610 AVDD.t588 AVDD.t587 AVDD.t588 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X611 AVDD.t586 AVDD.t585 AVDD.t586 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X612 AVSS.t129 AVSS.t128 AVSS.t129 AVSS.t77 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X613 AVDD IREF.t179 a_n13990_8177.t165 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X614 AVDD.t584 AVDD.t583 AVDD.t584 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X615 AVDD.t582 AVDD.t581 AVDD.t582 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X616 AVDD.t580 AVDD.t579 AVDD.t580 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X617 AVDD.t578 AVDD.t577 AVDD.t578 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X618 AVDD.t576 AVDD.t575 AVDD.t576 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X619 AVDD.t574 AVDD.t573 AVDD.t574 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X620 AVDD IREF.t180 a_n13990_8177.t164 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X621 AVDD.t572 AVDD.t571 AVDD.t572 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X622 AVDD a_5396_n6451.t207 a_5396_8177.t37 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X623 AVDD.t570 AVDD.t569 AVDD.t570 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X624 AVDD a_5396_n6451.t208 a_5396_9163.t36 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X625 AVDD.t568 AVDD.t567 AVDD.t568 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X626 VOUT a_n11317_n20927.t1 a_5396_9163.t101 AVDD.t121 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X627 AVDD.t566 AVDD.t565 AVDD.t566 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X628 AVDD.t564 AVDD.t563 AVDD.t564 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X629 AVDD IREF.t182 a_n13990_8177.t162 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X630 AVDD.t562 AVDD.t561 AVDD.t562 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X631 AVDD IREF.t185 a_n13990_8177.t159 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X632 AVDD a_5396_n6451.t209 a_5396_9163.t35 AVDD.t22 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X633 AVDD.t560 AVDD.t559 AVDD.t560 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X634 VOUT a_n11317_n20927.t1 a_5396_9163.t100 AVDD.t121 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X635 AVDD.t558 AVDD.t557 AVDD.t558 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X636 AVDD.t556 AVDD.t554 AVDD.t556 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X637 AVDD a_5396_n6451.t210 a_5396_8177.t36 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X638 AVDD.t553 AVDD.t552 AVDD.t553 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X639 AVDD.t551 AVDD.t550 AVDD.t551 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X640 AVDD.t549 AVDD.t548 AVDD.t549 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X641 AVDD a_5396_n6451.t211 a_5396_8177.t35 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X642 AVDD.t547 AVDD.t546 AVDD.t547 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X643 AVDD.t545 AVDD.t544 AVDD.t545 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X644 AVDD.t543 AVDD.t542 AVDD.t543 AVDD.t2 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X645 AVSS.t127 AVSS.t126 AVSS.t127 AVSS.t52 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X646 AVDD.t541 AVDD.t540 AVDD.t541 AVDD.t110 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X647 AVDD.t539 AVDD.t538 AVDD.t539 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X648 AVDD IREF.t16 IREF.t17 AVDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X649 AVDD.t537 AVDD.t536 AVDD.t537 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X650 AVDD.t535 AVDD.t534 AVDD.t535 AVDD.t110 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X651 AVDD.t533 AVDD.t532 AVDD.t533 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X652 AVDD.t531 AVDD.t530 AVDD.t531 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X653 AVSS.t125 AVSS.t124 AVSS.t125 AVSS.t46 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X654 AVSS a_n11737_n14973.t72 a_n13990_n6451.t46 AVSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X655 AVDD.t529 AVDD.t528 AVDD.t529 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X656 AVDD.t527 AVDD.t526 AVDD.t527 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X657 AVDD.t525 AVDD.t524 AVDD.t525 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X658 AVDD.t523 AVDD.t522 AVDD.t523 AVDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X659 AVDD.t521 AVDD.t520 AVDD.t521 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X660 AVDD.t519 AVDD.t518 AVDD.t519 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X661 AVDD IREF.t14 IREF.t15 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X662 AVDD IREF.t189 a_n13990_8177.t157 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X663 AVDD a_5396_n6451.t213 a_5396_8177.t33 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X664 AVDD.t517 AVDD.t516 AVDD.t517 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X665 AVDD.t515 AVDD.t514 AVDD.t515 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X666 AVDD.t513 AVDD.t512 AVDD.t513 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X667 AVDD.t511 AVDD.t510 AVDD.t511 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X668 AVDD.t509 AVDD.t508 AVDD.t509 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X669 AVDD.t507 AVDD.t506 AVDD.t507 AVDD.t92 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X670 AVDD.t505 AVDD.t504 AVDD.t505 AVDD.t110 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X671 AVDD.t503 AVDD.t502 AVDD.t503 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X672 AVDD.t501 AVDD.t500 AVDD.t501 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X673 AVDD a_5396_n6451.t215 a_5396_8177.t32 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X674 AVDD.t499 AVDD.t498 AVDD.t499 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X675 AVDD.t497 AVDD.t496 AVDD.t497 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X676 AVDD.t495 AVDD.t494 AVDD.t495 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X677 AVDD IREF.t191 a_n13990_8177.t155 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X678 AVDD IREF.t192 a_n13990_8177.t154 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X679 AVDD a_5396_n6451.t217 a_5396_8177.t31 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X680 AVDD IREF.t194 a_n11737_n15980.t10 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X681 AVDD.t493 AVDD.t492 AVDD.t493 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X682 AVSS.t123 AVSS.t122 AVSS.t123 AVSS.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X683 AVDD.t491 AVDD.t490 AVDD.t491 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X684 AVDD IREF.t195 a_n13990_8177.t152 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X685 AVDD.t489 AVDD.t488 AVDD.t489 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X686 AVDD a_5396_n6451.t218 a_5396_9163.t32 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X687 AVSS a_n11737_n14973.t77 a_n13990_n5465.t20 AVSS.t43 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X688 AVDD.t487 AVDD.t486 AVDD.t487 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X689 AVSS.t121 AVSS.t120 AVSS.t121 AVSS.t85 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X690 AVDD.t485 AVDD.t484 AVDD.t485 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X691 AVDD a_5396_n6451.t220 a_5396_9163.t31 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X692 AVDD.t483 AVDD.t482 AVDD.t483 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X693 AVDD IREF.t198 a_n13990_8177.t149 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X694 AVDD.t481 AVDD.t479 AVDD.t481 AVDD.t480 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X695 AVDD.t478 AVDD.t477 AVDD.t478 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X696 AVDD.t476 AVDD.t475 AVDD.t476 AVDD.t39 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X697 AVDD.t474 AVDD.t473 AVDD.t474 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X698 AVDD.t472 AVDD.t471 AVDD.t472 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X699 AVSS.t119 AVSS.t118 AVSS.t119 AVSS.t82 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X700 AVDD.t470 AVDD.t469 AVDD.t470 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X701 AVDD.t468 AVDD.t467 AVDD.t468 AVDD.t192 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X702 AVDD.t466 AVDD.t465 AVDD.t466 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X703 AVDD.t464 AVDD.t463 AVDD.t464 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X704 AVDD.t462 AVDD.t461 AVDD.t462 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X705 AVSS a_n11737_n14973.t78 a_n13990_n6451.t16 AVSS.t235 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X706 AVDD.t460 AVDD.t459 AVDD.t460 AVDD.t192 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X707 AVDD.t458 AVDD.t457 AVDD.t458 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X708 AVDD.t456 AVDD.t455 AVDD.t456 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X709 AVDD IREF.t201 a_n13990_8177.t147 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X710 AVDD IREF.t202 a_n13990_8177.t146 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X711 AVDD.t454 AVDD.t453 AVDD.t454 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X712 AVDD.t452 AVDD.t451 AVDD.t452 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X713 AVSS.t117 AVSS.t116 AVSS.t117 AVSS.t28 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X714 AVSS a_n11737_n14973.t79 a_n11317_n20927.t1 AVSS.t138 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X715 AVDD.t450 AVDD.t449 AVDD.t450 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X716 AVDD.t448 AVDD.t447 AVDD.t448 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X717 AVSS a_n11737_n14973.t80 a_n13990_n5465.t10 AVSS.t144 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X718 AVSS a_n11737_n14973.t81 a_n13990_n5465.t11 AVSS.t141 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X719 AVDD.t446 AVDD.t445 AVDD.t446 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X720 AVDD IREF.t203 a_n13990_8177.t145 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X721 AVDD.t444 AVDD.t443 AVDD.t444 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X722 AVDD a_5396_n6451.t223 a_5396_8177.t28 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X723 AVDD.t442 AVDD.t441 AVDD.t442 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X724 AVDD.t440 AVDD.t439 AVDD.t440 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X725 AVDD.t438 AVDD.t437 AVDD.t438 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X726 AVDD IREF.t204 a_n13990_8177.t144 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X727 AVDD.t436 AVDD.t435 AVDD.t436 AVDD.t2 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X728 VOUT a_n11317_n20927.t1 a_5396_9163.t99 AVDD.t110 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X729 VOUT a_n11737_n15980.t52 a_n13990_n5465.t33 AVSS.t1 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X730 VOUT a_n11737_n15980.t53 a_n13990_n5465.t32 AVSS.t2 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X731 AVDD.t434 AVDD.t433 AVDD.t434 AVDD.t177 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X732 AVDD.t432 AVDD.t431 AVDD.t432 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X733 AVSS.t115 AVSS.t113 AVSS.t115 AVSS.t114 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X734 AVDD.t430 AVDD.t429 AVDD.t430 AVDD.t195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X735 AVDD IREF.t205 a_n13990_8177.t143 AVDD.t252 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X736 AVSS a_n11737_n14973.t0 a_n11737_n14973.t1 AVSS.t133 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X737 AVDD a_5396_n6451.t224 a_5396_8177.t27 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X738 AVDD.t428 AVDD.t427 AVDD.t428 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X739 AVSS.t112 AVSS.t111 AVSS.t112 AVSS.t52 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X740 AVDD.t426 AVDD.t425 AVDD.t426 AVDD.t195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X741 AVDD IREF.t206 a_n13990_8177.t142 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X742 AVDD.t424 AVDD.t423 AVDD.t424 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X743 AVDD.t422 AVDD.t421 AVDD.t422 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X744 VOUT a_n11317_n20927.t7 a_5396_9163.t98 AVDD.t110 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X745 VOUT a_n11317_n20927.t1 a_5396_9163.t97 AVDD.t121 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X746 AVDD.t420 AVDD.t419 AVDD.t420 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X747 AVDD IREF.t209 a_n11737_n14973.t13 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X748 AVDD a_5396_n6451.t225 a_5396_9163.t29 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X749 AVDD.t418 AVDD.t417 AVDD.t418 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X750 AVDD.t416 AVDD.t415 AVDD.t416 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X751 AVDD a_5396_n6451.t226 a_5396_9163.t28 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X752 AVSS a_n11737_n14973.t86 a_n13990_n5465.t4 AVSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X753 AVDD.t414 AVDD.t413 AVDD.t414 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X754 AVDD.t412 AVDD.t411 AVDD.t412 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X755 VOUT a_n11737_n15980.t54 a_n13990_n5465.t31 AVSS.t16 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X756 VOUT a_n11317_n20927.t1 a_5396_9163.t96 AVDD.t121 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X757 AVDD IREF.t210 a_n11737_n14973.t12 AVDD.t810 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X758 VOUT a_n11737_n15980.t55 a_n13990_n5465.t30 AVSS.t13 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X759 AVDD.t410 AVDD.t409 AVDD.t410 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X760 AVDD IREF.t211 a_n13990_8177.t140 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X761 AVDD IREF.t212 a_n11737_n15980.t8 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X762 AVDD.t408 AVDD.t407 AVDD.t408 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X763 AVDD a_5396_n6451.t227 a_5396_8177.t26 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X764 AVDD a_5396_n6451.t229 a_5396_9163.t26 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X765 AVDD.t406 AVDD.t405 AVDD.t406 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X766 AVDD.t404 AVDD.t403 AVDD.t404 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X767 AVDD IREF.t213 a_n13990_8177.t139 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X768 AVSS.t110 AVSS.t109 AVSS.t110 AVSS.t99 nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X769 AVDD.t402 AVDD.t401 AVDD.t402 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X770 AVDD.t400 AVDD.t398 AVDD.t400 AVDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X771 AVDD.t397 AVDD.t396 AVDD.t397 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X772 AVDD.t395 AVDD.t393 AVDD.t395 AVDD.t394 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X773 AVDD.t392 AVDD.t391 AVDD.t392 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X774 AVSS a_n11737_n14973.t88 a_n13990_n5465.t17 AVSS.t222 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X775 AVDD.t390 AVDD.t389 AVDD.t390 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X776 AVDD.t388 AVDD.t387 AVDD.t388 AVDD.t13 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X777 AVDD.t386 AVDD.t385 AVDD.t386 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X778 AVDD IREF.t215 a_n13990_8177.t137 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X779 AVDD IREF.t216 a_n13990_8177.t136 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X780 AVDD.t384 AVDD.t383 AVDD.t384 AVDD.t155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X781 AVDD.t382 AVDD.t380 AVDD.t382 AVDD.t381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X782 AVDD.t379 AVDD.t377 AVDD.t379 AVDD.t378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X783 AVDD.t376 AVDD.t375 AVDD.t376 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X784 AVDD a_5396_n6451.t233 a_5396_9163.t25 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X785 AVDD a_5396_n6451.t234 a_5396_8177.t22 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X786 AVDD IREF.t219 a_n13990_8177.t134 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X787 AVDD.t374 AVDD.t372 AVDD.t374 AVDD.t373 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X788 AVSS.t108 AVSS.t107 AVSS.t108 AVSS.t77 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X789 VOUT a_n11317_n20927.t1 a_5396_9163.t95 AVDD.t200 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X790 AVDD.t371 AVDD.t370 AVDD.t371 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X791 AVDD.t369 AVDD.t368 AVDD.t369 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X792 AVDD.t367 AVDD.t365 AVDD.t367 AVDD.t366 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X793 AVSS.t106 AVSS.t105 AVSS.t106 AVSS.t55 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X794 AVDD.t364 AVDD.t363 AVDD.t364 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X795 AVDD.t362 AVDD.t361 AVDD.t362 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X796 AVSS.t104 AVSS.t103 AVSS.t104 AVSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X797 AVSS.t102 AVSS.t101 AVSS.t102 AVSS.t4 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X798 AVDD.t360 AVDD.t359 AVDD.t360 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X799 AVDD.t358 AVDD.t357 AVDD.t358 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X800 AVSS.t100 AVSS.t98 AVSS.t100 AVSS.t99 nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X801 AVDD IREF.t223 a_n13990_8177.t130 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X802 AVSS.t97 AVSS.t95 AVSS.t97 AVSS.t96 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X803 VOUT a_n11317_n20927.t1 a_5396_9163.t94 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X804 AVDD.t356 AVDD.t355 AVDD.t356 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X805 AVDD.t354 AVDD.t353 AVDD.t354 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X806 AVDD IREF.t224 a_n13990_8177.t129 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X807 AVDD a_5396_n6451.t236 a_5396_9163.t23 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X808 VOUT a_n11737_n15980.t58 a_n13990_n5465.t29 AVSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X809 AVSS.t94 AVSS.t93 AVSS.t94 AVSS.t46 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X810 AVDD.t352 AVDD.t351 AVDD.t352 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X811 AVDD a_5396_n6451.t237 a_5396_9163.t22 AVDD.t347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X812 AVDD a_5396_n6451.t238 a_5396_8177.t21 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X813 AVDD.t350 AVDD.t349 AVDD.t350 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X814 AVDD.t348 AVDD.t346 AVDD.t348 AVDD.t347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X815 AVDD.t345 AVDD.t344 AVDD.t345 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X816 AVDD IREF.t225 a_n13990_8177.t128 AVDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X817 AVDD.t343 AVDD.t342 AVDD.t343 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X818 AVDD.t341 AVDD.t340 AVDD.t341 AVDD.t195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X819 AVDD.t339 AVDD.t337 AVDD.t339 AVDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X820 AVDD.t336 AVDD.t334 AVDD.t336 AVDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X821 AVDD.t333 AVDD.t332 AVDD.t333 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X822 AVSS.t92 AVSS.t91 AVSS.t92 AVSS.t37 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X823 IREF IREF.t12 AVDD.t1705 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X824 AVSS a_n11737_n14973.t91 a_n13990_n6451.t21 AVSS.t201 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X825 AVDD.t331 AVDD.t330 AVDD.t331 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X826 AVDD.t329 AVDD.t327 AVDD.t329 AVDD.t328 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X827 AVDD.t326 AVDD.t325 AVDD.t326 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X828 IREF IREF.t10 AVDD.t1704 AVDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X829 AVDD.t324 AVDD.t322 AVDD.t324 AVDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X830 AVDD a_5396_n6451.t243 a_5396_8177.t19 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X831 AVDD.t321 AVDD.t320 AVDD.t321 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X832 AVDD.t319 AVDD.t318 AVDD.t319 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X833 AVDD.t317 AVDD.t316 AVDD.t317 AVDD.t155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X834 AVDD.t315 AVDD.t314 AVDD.t315 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X835 AVDD.t313 AVDD.t312 AVDD.t313 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X836 AVDD a_5396_n6451.t244 a_5396_9163.t18 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X837 AVDD.t311 AVDD.t310 AVDD.t311 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X838 AVDD.t309 AVDD.t308 AVDD.t309 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X839 AVDD a_5396_n6451.t246 a_5396_9163.t16 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X840 AVSS.t90 AVSS.t89 AVSS.t90 AVSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X841 AVSS.t88 AVSS.t87 AVSS.t88 AVSS.t2 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X842 AVSS.t86 AVSS.t84 AVSS.t86 AVSS.t85 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X843 AVDD a_5396_n6451.t247 a_5396_8177.t18 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X844 AVDD.t307 AVDD.t306 AVDD.t307 AVDD.t192 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X845 AVSS a_n11737_n14973.t92 a_n13990_n5465.t25 AVSS.t235 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X846 AVDD.t305 AVDD.t304 AVDD.t305 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X847 AVDD IREF.t233 a_n13990_8177.t122 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X848 AVDD.t303 AVDD.t302 AVDD.t303 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X849 AVSS.t83 AVSS.t81 AVSS.t83 AVSS.t82 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X850 AVDD a_5396_n6451.t248 a_5396_9163.t15 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X851 AVDD.t301 AVDD.t300 AVDD.t301 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X852 AVDD.t299 AVDD.t298 AVDD.t299 AVDD.t155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X853 AVSS.t80 AVSS.t79 AVSS.t80 AVSS.t28 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X854 AVDD.t297 AVDD.t296 AVDD.t297 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X855 AVDD.t295 AVDD.t293 AVDD.t295 AVDD.t294 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X856 AVSS.t78 AVSS.t76 AVSS.t78 AVSS.t77 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X857 AVDD.t292 AVDD.t290 AVDD.t292 AVDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X858 AVDD IREF.t236 a_n13990_8177.t119 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X859 AVDD.t289 AVDD.t288 AVDD.t289 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X860 AVDD a_5396_n6451.t251 a_5396_9163.t13 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X861 AVDD a_5396_n6451.t252 a_5396_8177.t16 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X862 AVDD a_5396_n6451.t253 a_5396_9163.t12 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X863 AVDD.t287 AVDD.t286 AVDD.t287 AVDD.t152 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X864 AVDD.t285 AVDD.t284 AVDD.t285 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X865 AVDD.t283 AVDD.t281 AVDD.t283 AVDD.t282 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X866 AVDD.t280 AVDD.t278 AVDD.t280 AVDD.t279 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X867 AVDD.t277 AVDD.t276 AVDD.t277 AVDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X868 AVSS.t75 AVSS.t74 AVSS.t75 AVSS.t49 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X869 AVDD IREF.t8 IREF.t9 AVDD.t810 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X870 AVDD.t275 AVDD.t274 AVDD.t275 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X871 AVDD.t273 AVDD.t272 AVDD.t273 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X872 AVDD IREF.t6 IREF.t7 AVDD.t638 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X873 AVDD.t271 AVDD.t270 AVDD.t271 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X874 AVDD.t269 AVDD.t268 AVDD.t269 AVDD.t135 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X875 AVDD.t267 AVDD.t266 AVDD.t267 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X876 AVDD.t265 AVDD.t263 AVDD.t265 AVDD.t264 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X877 AVDD.t262 AVDD.t261 AVDD.t262 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X878 AVDD.t260 AVDD.t259 AVDD.t260 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X879 AVDD.t258 AVDD.t257 AVDD.t258 AVDD.t92 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X880 AVDD.t256 AVDD.t254 AVDD.t256 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X881 AVDD.t253 AVDD.t251 AVDD.t253 AVDD.t252 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X882 AVSS.t73 AVSS.t72 AVSS.t73 AVSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X883 AVSS.t71 AVSS.t69 AVSS.t71 AVSS.t70 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X884 AVDD.t250 AVDD.t249 AVDD.t250 AVDD.t177 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X885 AVSS.t68 AVSS.t66 AVSS.t68 AVSS.t67 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X886 AVDD.t248 AVDD.t247 AVDD.t248 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X887 AVDD IREF.t240 a_n13990_8177.t116 AVDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X888 AVDD.t246 AVDD.t245 AVDD.t246 AVDD.t180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X889 AVDD.t244 AVDD.t243 AVDD.t244 AVDD.t177 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X890 AVDD.t242 AVDD.t240 AVDD.t242 AVDD.t241 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X891 AVDD.t239 AVDD.t237 AVDD.t239 AVDD.t238 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X892 AVDD.t236 AVDD.t235 AVDD.t236 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X893 AVDD.t234 AVDD.t232 AVDD.t234 AVDD.t233 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X894 AVSS.t65 AVSS.t64 AVSS.t65 AVSS.t4 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X895 AVSS.t63 AVSS.t62 AVSS.t63 AVSS.t37 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X896 AVDD a_5396_n6451.t257 a_5396_9163.t10 AVDD.t226 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X897 AVDD.t231 AVDD.t230 AVDD.t231 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X898 AVDD.t229 AVDD.t228 AVDD.t229 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X899 AVDD.t227 AVDD.t225 AVDD.t227 AVDD.t226 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X900 AVDD.t224 AVDD.t223 AVDD.t224 AVDD.t121 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X901 AVDD.t222 AVDD.t221 AVDD.t222 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X902 AVDD.t220 AVDD.t219 AVDD.t220 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X903 AVDD IREF.t242 a_n11737_n15980.t5 AVDD.t282 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X904 AVDD.t218 AVDD.t217 AVDD.t218 AVDD.t192 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X905 AVDD.t216 AVDD.t215 AVDD.t216 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X906 VOUT a_n11317_n20927.t1 a_5396_9163.t93 AVDD.t381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X907 AVSS a_n11737_n14973.t96 a_n13990_n6451.t8 AVSS.t222 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X908 AVSS.t61 AVSS.t60 AVSS.t61 AVSS.t31 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X909 AVDD IREF.t243 a_n11737_n15980.t4 AVDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X910 AVDD.t214 AVDD.t213 AVDD.t214 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X911 AVDD.t212 AVDD.t211 AVDD.t212 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X912 a_n5579_n20820# a_n11737_n15980.t63 a_n6139_n20267# AVSS.t99 nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X913 AVDD.t210 AVDD.t209 AVDD.t210 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X914 AVDD.t208 AVDD.t207 AVDD.t208 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X915 AVDD.t206 AVDD.t204 AVDD.t206 AVDD.t205 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X916 AVDD.t203 AVDD.t202 AVDD.t203 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X917 a_n1533_n16909# a_n11317_n20927.t1 a_n2101_n16909# AVDD.t394 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X918 AVDD.t201 AVDD.t199 AVDD.t201 AVDD.t200 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X919 AVDD IREF.t244 a_n13990_8177.t114 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X920 AVDD IREF.t246 a_n13990_8177.t112 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X921 AVDD.t198 AVDD.t197 AVDD.t198 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X922 AVDD.t196 AVDD.t194 AVDD.t196 AVDD.t195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X923 AVDD.t193 AVDD.t191 AVDD.t193 AVDD.t192 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X924 AVDD.t190 AVDD.t189 AVDD.t190 AVDD.t130 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X925 AVDD.t188 AVDD.t187 AVDD.t188 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X926 AVDD.t186 AVDD.t184 AVDD.t186 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X927 AVDD.t183 AVDD.t182 AVDD.t183 AVDD.t152 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X928 AVDD.t181 AVDD.t179 AVDD.t181 AVDD.t180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X929 AVSS.t59 AVSS.t57 AVSS.t59 AVSS.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X930 VOUT a_n11317_n20927.t1 a_5396_9163.t92 AVDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X931 VOUT a_n11737_n15980.t64 a_n13990_n5465.t28 AVSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X932 AVDD a_5396_n6451.t264 a_5396_9163.t8 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X933 AVDD.t178 AVDD.t176 AVDD.t178 AVDD.t177 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X934 AVSS.t56 AVSS.t54 AVSS.t56 AVSS.t55 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X935 AVDD.t175 AVDD.t173 AVDD.t175 AVDD.t174 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X936 AVDD.t172 AVDD.t171 AVDD.t172 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X937 AVDD a_5396_n6451.t265 a_5396_8177.t8 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X938 AVDD.t170 AVDD.t169 AVDD.t170 AVDD.t135 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X939 AVDD.t168 AVDD.t167 AVDD.t168 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X940 AVDD.t166 AVDD.t165 AVDD.t166 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X941 VOUT a_n11317_n20927.t1 a_5396_9163.t91 AVDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X942 AVSS.t53 AVSS.t51 AVSS.t53 AVSS.t52 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X943 AVDD.t164 AVDD.t163 AVDD.t164 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X944 AVDD.t162 AVDD.t161 AVDD.t162 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X945 AVDD.t160 AVDD.t159 AVDD.t160 AVDD.t155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X946 AVDD.t158 AVDD.t157 AVDD.t158 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X947 AVDD IREF.t250 a_n11737_n15980.t3 AVDD.t717 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X948 AVDD.t156 AVDD.t154 AVDD.t156 AVDD.t155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X949 AVDD.t153 AVDD.t151 AVDD.t153 AVDD.t152 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X950 AVDD.t150 AVDD.t149 AVDD.t150 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X951 AVDD.t148 AVDD.t146 AVDD.t148 AVDD.t147 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X952 AVDD IREF.t251 a_n13990_8177.t108 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X953 AVDD.t145 AVDD.t144 AVDD.t145 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X954 AVDD.t143 AVDD.t142 AVDD.t143 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X955 AVDD IREF.t252 a_n11737_n14973.t11 AVDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X956 AVDD.t141 AVDD.t139 AVDD.t141 AVDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X957 AVDD.t138 AVDD.t137 AVDD.t138 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X958 IREF IREF.t4 AVDD.t1798 AVDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X959 AVDD.t136 AVDD.t134 AVDD.t136 AVDD.t135 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X960 AVSS a_n11737_n14973.t101 a_n13990_n5465.t0 AVSS.t201 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X961 AVDD.t133 AVDD.t132 AVDD.t133 AVDD.t121 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X962 AVDD.t131 AVDD.t129 AVDD.t131 AVDD.t130 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X963 AVSS.t50 AVSS.t48 AVSS.t50 AVSS.t49 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X964 AVDD.t128 AVDD.t127 AVDD.t128 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X965 AVSS.t47 AVSS.t45 AVSS.t47 AVSS.t46 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X966 AVSS a_n11737_n14973.t102 a_n13990_n5465.t1 AVSS.t114 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X967 a_n2101_n16909# a_n11317_n20927.t1 a_n2631_n17634# AVDD.t328 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X968 AVSS.t44 AVSS.t42 AVSS.t44 AVSS.t43 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X969 AVDD IREF.t255 a_n13990_8177.t106 AVDD.t152 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X970 AVDD.t126 AVDD.t125 AVDD.t126 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X971 AVDD.t124 AVDD.t123 AVDD.t124 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X972 AVDD.t122 AVDD.t120 AVDD.t122 AVDD.t121 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X973 AVDD.t119 AVDD.t117 AVDD.t119 AVDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X974 AVDD IREF.t256 a_n13990_8177.t105 AVDD.t255 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X975 AVDD.t116 AVDD.t115 AVDD.t116 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X976 AVDD.t114 AVDD.t112 AVDD.t114 AVDD.t113 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X977 AVDD IREF.t2 IREF.t3 AVDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X978 AVSS.t41 AVSS.t39 AVSS.t41 AVSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X979 AVDD.t111 AVDD.t109 AVDD.t111 AVDD.t110 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X980 AVDD.t108 AVDD.t107 AVDD.t108 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X981 AVDD.t106 AVDD.t105 AVDD.t106 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X982 AVDD.t104 AVDD.t103 AVDD.t104 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X983 AVDD.t102 AVDD.t101 AVDD.t102 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X984 AVDD IREF.t258 a_n13990_8177.t103 AVDD.t233 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X985 AVDD.t100 AVDD.t99 AVDD.t100 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X986 AVDD.t98 AVDD.t96 AVDD.t98 AVDD.t97 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X987 AVDD.t95 AVDD.t94 AVDD.t95 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X988 AVDD.t93 AVDD.t91 AVDD.t93 AVDD.t92 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X989 AVDD.t90 AVDD.t89 AVDD.t90 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X990 AVDD.t88 AVDD.t86 AVDD.t88 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X991 AVDD.t85 AVDD.t84 AVDD.t85 AVDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X992 AVDD.t83 AVDD.t81 AVDD.t83 AVDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X993 AVDD.t80 AVDD.t78 AVDD.t80 AVDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X994 AVDD.t77 AVDD.t76 AVDD.t77 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X995 AVDD.t75 AVDD.t74 AVDD.t75 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X996 AVDD a_5396_n6451.t272 a_5396_8177.t4 AVDD.t241 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X997 AVDD.t73 AVDD.t72 AVDD.t73 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X998 AVSS.t38 AVSS.t36 AVSS.t38 AVSS.t37 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X999 AVDD.t71 AVDD.t69 AVDD.t71 AVDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1000 AVDD.t68 AVDD.t66 AVDD.t68 AVDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1001 AVDD IREF.t0 IREF.t1 AVDD.t810 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1002 AVDD IREF.t264 a_n13990_8177.t100 AVDD.t33 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1003 AVSS.t35 AVSS.t33 AVSS.t35 AVSS.t34 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X1004 AVSS.t32 AVSS.t30 AVSS.t32 AVSS.t31 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1005 AVDD.t65 AVDD.t64 AVDD.t65 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1006 AVDD.t63 AVDD.t61 AVDD.t63 AVDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1007 AVDD.t60 AVDD.t58 AVDD.t60 AVDD.t59 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1008 AVDD.t57 AVDD.t55 AVDD.t57 AVDD.t56 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1009 AVDD.t54 AVDD.t52 AVDD.t54 AVDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1010 AVDD a_5396_n6451.t274 a_5396_9163.t3 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1011 AVDD.t51 AVDD.t50 AVDD.t51 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1012 AVDD.t49 AVDD.t48 AVDD.t49 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1013 AVSS.t29 AVSS.t27 AVSS.t29 AVSS.t28 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1014 VOUT a_n11317_n20927.t1 a_5396_9163.t90 AVDD.t59 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1015 AVSS.t26 AVSS.t24 AVSS.t26 AVSS.t25 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1016 AVSS.t23 AVSS.t21 AVSS.t23 AVSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1017 AVSS.t20 AVSS.t18 AVSS.t20 AVSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1018 AVSS.t17 AVSS.t15 AVSS.t17 AVSS.t16 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1019 AVDD.t47 AVDD.t46 AVDD.t47 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1020 AVSS.t14 AVSS.t12 AVSS.t14 AVSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1021 AVDD.t45 AVDD.t43 AVDD.t45 AVDD.t44 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1022 VOUT a_n11317_n20927.t1 a_5396_9163.t89 AVDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1023 AVDD.t42 AVDD.t41 AVDD.t42 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1024 AVDD.t40 AVDD.t38 AVDD.t40 AVDD.t39 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1025 AVDD.t37 AVDD.t35 AVDD.t37 AVDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1026 AVDD.t34 AVDD.t32 AVDD.t34 AVDD.t33 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1027 AVSS.t11 AVSS.t9 AVSS.t11 AVSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1028 AVDD IREF.t270 a_n13990_8177.t94 AVDD.t185 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1029 AVSS.t8 AVSS.t6 AVSS.t8 AVSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1030 AVDD.t31 AVDD.t29 AVDD.t31 AVDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1031 AVDD.t28 AVDD.t26 AVDD.t28 AVDD.t27 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1032 AVDD.t25 AVDD.t24 AVDD.t25 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1033 AVDD.t23 AVDD.t21 AVDD.t23 AVDD.t22 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1034 AVDD.t20 AVDD.t18 AVDD.t20 AVDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1035 VOUT a_n11317_n20927.t1 a_5396_9163.t88 AVDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1036 AVDD.t17 AVDD.t15 AVDD.t17 AVDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1037 AVDD.t14 AVDD.t12 AVDD.t14 AVDD.t13 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1038 AVDD.t11 AVDD.t10 AVDD.t11 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1039 AVSS.t5 AVSS.t3 AVSS.t5 AVSS.t4 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1040 AVDD.t9 AVDD.t7 AVDD.t9 AVDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1041 AVDD.t6 AVDD.t4 AVDD.t6 AVDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1042 AVDD a_5396_n6451.t280 a_5396_8177.t1 AVDD.t87 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1043 AVDD.t3 AVDD.t1 AVDD.t3 AVDD.t2 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
R0 AVDD.n1124 AVDD.n954 714.056
R1 AVDD.n1124 AVDD.n953 712.232
R2 AVDD.n1129 AVDD.n954 707.59
R3 AVDD.n1129 AVDD.n953 705.766
R4 AVDD.n1305 AVDD.n41 647.574
R5 AVDD.n2146 AVDD.n4 647.574
R6 AVDD.n1482 AVDD.n1 647.574
R7 AVDD.n93 AVDD.n92 647.574
R8 AVDD.n23 AVDD.n21 647.574
R9 AVDD.n1451 AVDD.n113 647.574
R10 AVDD.n100 AVDD.n94 647.574
R11 AVDD.n1307 AVDD.n707 647.574
R12 AVDD.n883 AVDD.n9 647.574
R13 AVDD.n119 AVDD.n11 647.574
R14 AVDD.n493 AVDD.n95 647.574
R15 AVDD.n1241 AVDD.n710 647.574
R16 AVDD.n2181 AVDD.n20 647.574
R17 AVDD.n120 AVDD.n14 647.574
R18 AVDD.n561 AVDD.n96 647.574
R19 AVDD.n708 AVDD.n36 647.574
R20 AVDD.n2153 AVDD.n41 642.269
R21 AVDD.n2220 AVDD.n4 642.269
R22 AVDD.n1495 AVDD.n1482 642.269
R23 AVDD.n93 AVDD.n91 642.269
R24 AVDD.n21 AVDD.n6 642.269
R25 AVDD.n1497 AVDD.n113 642.269
R26 AVDD.n99 AVDD.n94 642.269
R27 AVDD.n707 AVDD.n39 642.269
R28 AVDD.n2218 AVDD.n9 642.269
R29 AVDD.n119 AVDD.n116 642.269
R30 AVDD.n608 AVDD.n95 642.269
R31 AVDD.n710 AVDD.n38 642.269
R32 AVDD.n2181 AVDD.n7 642.269
R33 AVDD.n120 AVDD.n115 642.269
R34 AVDD.n606 AVDD.n96 642.269
R35 AVDD.n2155 AVDD.n36 642.269
R36 AVDD.n1305 AVDD.n40 640.197
R37 AVDD.n2146 AVDD.n3 640.197
R38 AVDD.n117 AVDD.n1 640.197
R39 AVDD.n1523 AVDD.n92 640.197
R40 AVDD.n2179 AVDD.n23 640.197
R41 AVDD.n1451 AVDD.n112 640.197
R42 AVDD.n1521 AVDD.n100 640.197
R43 AVDD.n1307 AVDD.n696 640.197
R44 AVDD.n883 AVDD.n8 640.197
R45 AVDD.n1480 AVDD.n11 640.197
R46 AVDD.n493 AVDD.n98 640.197
R47 AVDD.n1241 AVDD.n709 640.197
R48 AVDD.n22 AVDD.n20 640.197
R49 AVDD.n121 AVDD.n14 640.197
R50 AVDD.n561 AVDD.n97 640.197
R51 AVDD.n708 AVDD.n35 640.197
R52 AVDD.n2153 AVDD.n40 634.891
R53 AVDD.n2220 AVDD.n3 634.891
R54 AVDD.n1495 AVDD.n117 634.891
R55 AVDD.n1523 AVDD.n91 634.891
R56 AVDD.n2179 AVDD.n6 634.891
R57 AVDD.n1497 AVDD.n112 634.891
R58 AVDD.n1521 AVDD.n99 634.891
R59 AVDD.n696 AVDD.n39 634.891
R60 AVDD.n2218 AVDD.n8 634.891
R61 AVDD.n1480 AVDD.n116 634.891
R62 AVDD.n608 AVDD.n98 634.891
R63 AVDD.n709 AVDD.n38 634.891
R64 AVDD.n22 AVDD.n7 634.891
R65 AVDD.n121 AVDD.n115 634.891
R66 AVDD.n606 AVDD.n97 634.891
R67 AVDD.n2155 AVDD.n35 634.891
R68 AVDD.n1049 AVDD.n956 351.805
R69 AVDD.n1122 AVDD.n956 351.639
R70 AVDD.n1049 AVDD.n955 350.479
R71 AVDD.n1122 AVDD.n955 350.313
R72 AVDD.n407 AVDD.n148 322.38
R73 AVDD.n604 AVDD.n409 289.171
R74 AVDD.n368 AVDD.n149 289.171
R75 AVDD.n402 AVDD.n149 267.75
R76 AVDD.n409 AVDD.n407 255.06
R77 AVDD.n402 AVDD.n148 255.06
R78 AVDD.t328 AVDD.t13 85.1494
R79 AVDD.t130 AVDD.t39 85.1494
R80 AVDD.t810 AVDD.t180 85.1494
R81 AVDD.t373 AVDD.t2 81.7244
R82 AVDD.t638 AVDD.t875 79.7265
R83 AVDD.t2 AVDD.t264 79.5362
R84 AVDD.n1127 AVDD.t27 68.5002
R85 AVDD.t394 AVDD.t328 54.0391
R86 AVDD.t39 AVDD.t555 54.0391
R87 AVDD.t555 AVDD.t480 54.0391
R88 AVDD.t480 AVDD.t282 54.0391
R89 AVDD.t717 AVDD.t638 54.0391
R90 AVDD.t875 AVDD.t366 54.0391
R91 AVDD.t366 AVDD.t323 54.0391
R92 AVDD.t323 AVDD.t810 54.0391
R93 AVDD.t27 AVDD.n1125 50.3287
R94 AVDD.n2219 AVDD.n5 46.8594
R95 AVDD.n1049 AVDD.t373 45.4522
R96 AVDD.t180 AVDD.n1124 45.3596
R97 AVDD.n1123 AVDD.t13 45.2864
R98 AVDD.n1128 AVDD.t130 45.2864
R99 AVDD.n1048 AVDD.t394 37.9607
R100 AVDD.t67 AVDD.t44 31.8205
R101 AVDD.t79 AVDD.t241 31.8205
R102 AVDD.t177 AVDD.t56 31.8205
R103 AVDD.t22 AVDD.t113 31.8205
R104 AVDD.t294 AVDD.t70 31.8205
R105 AVDD.t16 AVDD.t335 31.8205
R106 AVDD.t33 AVDD.t62 31.8205
R107 AVDD.t347 AVDD.t381 29.7939
R108 AVDD.t192 AVDD.t59 29.7939
R109 AVDD.t200 AVDD.t226 29.7939
R110 AVDD.t155 AVDD.t338 29.7939
R111 AVDD.t5 AVDD.t152 29.7939
R112 AVDD.t195 AVDD.t252 29.7939
R113 AVDD.t82 AVDD.t238 29.7939
R114 AVDD.t233 AVDD.t92 29.7939
R115 AVDD.t44 AVDD.t19 20.1946
R116 AVDD.t19 AVDD.t121 20.1946
R117 AVDD.t121 AVDD.t347 20.1946
R118 AVDD.t59 AVDD.t87 20.1946
R119 AVDD.t279 AVDD.t192 20.1946
R120 AVDD.t291 AVDD.t279 20.1946
R121 AVDD.t241 AVDD.t291 20.1946
R122 AVDD.t147 AVDD.t177 20.1946
R123 AVDD.t110 AVDD.t147 20.1946
R124 AVDD.t226 AVDD.t110 20.1946
R125 AVDD.t174 AVDD.t155 20.1946
R126 AVDD.t338 AVDD.t399 20.1946
R127 AVDD.t399 AVDD.t118 20.1946
R128 AVDD.t118 AVDD.t22 20.1946
R129 AVDD.t140 AVDD.t294 20.1946
R130 AVDD.t135 AVDD.t140 20.1946
R131 AVDD.t152 AVDD.t135 20.1946
R132 AVDD.t252 AVDD.t97 20.1946
R133 AVDD.t53 AVDD.t195 20.1946
R134 AVDD.t30 AVDD.t53 20.1946
R135 AVDD.t335 AVDD.t30 20.1946
R136 AVDD.t205 AVDD.t255 20.1946
R137 AVDD.t255 AVDD.t36 20.1946
R138 AVDD.t36 AVDD.t82 20.1946
R139 AVDD.t185 AVDD.t233 20.1946
R140 AVDD.t92 AVDD.t378 20.1946
R141 AVDD.t378 AVDD.t0 20.1946
R142 AVDD.t0 AVDD.t33 20.1946
R143 AVDD.n1522 AVDD.t381 19.0569
R144 AVDD.n1481 AVDD.t200 19.0569
R145 AVDD.n2180 AVDD.t5 19.0569
R146 AVDD.t238 AVDD.n1126 19.0569
R147 AVDD.n607 AVDD.t67 16.9237
R148 AVDD.n114 AVDD.t79 16.9237
R149 AVDD.n1496 AVDD.t56 16.9237
R150 AVDD.t113 AVDD.n5 16.9237
R151 AVDD.n2219 AVDD.t70 16.9237
R152 AVDD.n37 AVDD.t16 16.9237
R153 AVDD.n2154 AVDD.t8 16.9237
R154 AVDD.n1306 AVDD.t62 16.9237
R155 AVDD.n1127 AVDD.t8 16.4971
R156 AVDD.t264 AVDD.n1048 16.0789
R157 AVDD.n1127 AVDD.t205 15.3239
R158 AVDD.n1128 AVDD.n1123 13.7004
R159 AVDD.t282 AVDD.n1127 11.2268
R160 AVDD.n0 AVDD.t431 8.10567
R161 AVDD.n2224 AVDD.t953 8.10567
R162 AVDD.n2223 AVDD.t854 8.10567
R163 AVDD.n1439 AVDD.t923 8.10567
R164 AVDD.n1440 AVDD.t1105 8.10567
R165 AVDD.n1442 AVDD.t349 8.10567
R166 AVDD.n0 AVDD.t1187 8.10567
R167 AVDD.n2224 AVDD.t415 8.10567
R168 AVDD.n2223 AVDD.t320 8.10567
R169 AVDD.n1439 AVDD.t391 8.10567
R170 AVDD.n1440 AVDD.t587 8.10567
R171 AVDD.n1442 AVDD.t1083 8.10567
R172 AVDD.n1446 AVDD.t981 8.10567
R173 AVDD.n1448 AVDD.t207 8.10567
R174 AVDD.n1449 AVDD.t69 8.10567
R175 AVDD.n1454 AVDD.t211 8.10567
R176 AVDD.n1455 AVDD.t72 8.10567
R177 AVDD.n1457 AVDD.t676 8.10567
R178 AVDD.n1446 AVDD.t441 8.10567
R179 AVDD.n1448 AVDD.t959 8.10567
R180 AVDD.n1449 AVDD.t866 8.10567
R181 AVDD.n1454 AVDD.t221 8.10567
R182 AVDD.n1455 AVDD.t112 8.10567
R183 AVDD.n1457 AVDD.t694 8.10567
R184 AVDD.n1462 AVDD.t680 8.10567
R185 AVDD.n1460 AVDD.t1177 8.10567
R186 AVDD.n1459 AVDD.t1059 8.10567
R187 AVDD.n2215 AVDD.t1065 8.10567
R188 AVDD.n2214 AVDD.t759 8.10567
R189 AVDD.n2212 AVDD.t848 8.10567
R190 AVDD.n1462 AVDD.t702 8.10567
R191 AVDD.n1460 AVDD.t1191 8.10567
R192 AVDD.n1459 AVDD.t1069 8.10567
R193 AVDD.n2215 AVDD.t1089 8.10567
R194 AVDD.n2214 AVDD.t261 8.10567
R195 AVDD.n2212 AVDD.t314 8.10567
R196 AVDD.n2208 AVDD.t1225 8.10567
R197 AVDD.n2206 AVDD.t668 8.10567
R198 AVDD.n2205 AVDD.t793 8.10567
R199 AVDD.n2201 AVDD.t781 8.10567
R200 AVDD.n2200 AVDD.t889 8.10567
R201 AVDD.n2198 AVDD.t370 8.10567
R202 AVDD.n2208 AVDD.t725 8.10567
R203 AVDD.n2206 AVDD.t127 8.10567
R204 AVDD.n2205 AVDD.t266 8.10567
R205 AVDD.n2201 AVDD.t247 8.10567
R206 AVDD.n2200 AVDD.t353 8.10567
R207 AVDD.n2198 AVDD.t1119 8.10567
R208 AVDD.n72 AVDD.t137 8.10567
R209 AVDD.n71 AVDD.t1007 8.10567
R210 AVDD.n164 AVDD.t1263 8.10567
R211 AVDD.n161 AVDD.t421 8.10567
R212 AVDD.n160 AVDD.t383 8.10567
R213 AVDD.n171 AVDD.t670 8.10567
R214 AVDD.n159 AVDD.t1075 8.10567
R215 AVDD.n158 AVDD.t1107 8.10567
R216 AVDD.n179 AVDD.t109 8.10567
R217 AVDD.n156 AVDD.t652 8.10567
R218 AVDD.n155 AVDD.t933 8.10567
R219 AVDD.n45 AVDD.t1207 8.10567
R220 AVDD.n44 AVDD.t947 8.10567
R221 AVDD.n1737 AVDD.t52 8.10567
R222 AVDD.n1734 AVDD.t1063 8.10567
R223 AVDD.n1733 AVDD.t1135 8.10567
R224 AVDD.n1744 AVDD.t712 8.10567
R225 AVDD.n1732 AVDD.t417 8.10567
R226 AVDD.n1731 AVDD.t286 8.10567
R227 AVDD.n1752 AVDD.t268 8.10567
R228 AVDD.n69 AVDD.t642 8.10567
R229 AVDD.n68 AVDD.t1167 8.10567
R230 AVDD.n2141 AVDD.t46 8.10567
R231 AVDD.n2143 AVDD.t583 8.10567
R232 AVDD.n2144 AVDD.t451 8.10567
R233 AVDD.n2150 AVDD.t550 8.10567
R234 AVDD.n2149 AVDD.t751 8.10567
R235 AVDD.n2147 AVDD.t1235 8.10567
R236 AVDD.n2141 AVDD.t167 8.10567
R237 AVDD.n2143 AVDD.t690 8.10567
R238 AVDD.n2144 AVDD.t577 8.10567
R239 AVDD.n2150 AVDD.t650 8.10567
R240 AVDD.n2149 AVDD.t862 8.10567
R241 AVDD.n2147 AVDD.t48 8.10567
R242 AVDD.n2161 AVDD.t605 8.10567
R243 AVDD.n2159 AVDD.t1099 8.10567
R244 AVDD.n2158 AVDD.t999 8.10567
R245 AVDD.n1346 AVDD.t881 8.10567
R246 AVDD.n1347 AVDD.t773 8.10567
R247 AVDD.n2161 AVDD.t719 8.10567
R248 AVDD.n2159 AVDD.t1205 8.10567
R249 AVDD.n2158 AVDD.t1095 8.10567
R250 AVDD.n1346 AVDD.t457 8.10567
R251 AVDD.n1347 AVDD.t357 8.10567
R252 AVDD.n704 AVDD.t103 8.10567
R253 AVDD.n1317 AVDD.t664 8.10567
R254 AVDD.n702 AVDD.t284 8.10567
R255 AVDD.n1322 AVDD.t965 8.10567
R256 AVDD.n699 AVDD.t903 8.10567
R257 AVDD.n698 AVDD.t526 8.10567
R258 AVDD.n1329 AVDD.t905 8.10567
R259 AVDD.n694 AVDD.t500 8.10567
R260 AVDD.n1335 AVDD.t89 8.10567
R261 AVDD.n692 AVDD.t471 8.10567
R262 AVDD.n1340 AVDD.t747 8.10567
R263 AVDD.n689 AVDD.t1097 8.10567
R264 AVDD.n688 AVDD.t7 8.10567
R265 AVDD.n686 AVDD.t937 8.10567
R266 AVDD.n1353 AVDD.t1157 8.10567
R267 AVDD.n684 AVDD.t1067 8.10567
R268 AVDD.n1358 AVDD.t494 8.10567
R269 AVDD.n681 AVDD.t425 8.10567
R270 AVDD.n680 AVDD.t1015 8.10567
R271 AVDD.n1365 AVDD.t96 8.10567
R272 AVDD.n677 AVDD.t4 8.10567
R273 AVDD.n1371 AVDD.t593 8.10567
R274 AVDD.n675 AVDD.t1035 8.10567
R275 AVDD.n1376 AVDD.t1125 8.10567
R276 AVDD.n672 AVDD.t1209 8.10567
R277 AVDD.n704 AVDD.t115 8.10567
R278 AVDD.n1317 AVDD.t672 8.10567
R279 AVDD.n702 AVDD.t288 8.10567
R280 AVDD.n1322 AVDD.t971 8.10567
R281 AVDD.n699 AVDD.t909 8.10567
R282 AVDD.n698 AVDD.t532 8.10567
R283 AVDD.n1329 AVDD.t911 8.10567
R284 AVDD.n694 AVDD.t508 8.10567
R285 AVDD.n1335 AVDD.t101 8.10567
R286 AVDD.n692 AVDD.t484 8.10567
R287 AVDD.n1340 AVDD.t755 8.10567
R288 AVDD.n689 AVDD.t1103 8.10567
R289 AVDD.n688 AVDD.t24 8.10567
R290 AVDD.n686 AVDD.t941 8.10567
R291 AVDD.n1353 AVDD.t1165 8.10567
R292 AVDD.n684 AVDD.t1081 8.10567
R293 AVDD.n1358 AVDD.t502 8.10567
R294 AVDD.n681 AVDD.t429 8.10567
R295 AVDD.n680 AVDD.t1019 8.10567
R296 AVDD.n1365 AVDD.t105 8.10567
R297 AVDD.n677 AVDD.t10 8.10567
R298 AVDD.n1371 AVDD.t599 8.10567
R299 AVDD.n675 AVDD.t1045 8.10567
R300 AVDD.n1376 AVDD.t1133 8.10567
R301 AVDD.n672 AVDD.t1215 8.10567
R302 AVDD.n1311 AVDD.t625 8.10567
R303 AVDD.n1310 AVDD.t514 8.10567
R304 AVDD.n805 AVDD.t520 8.10567
R305 AVDD.n806 AVDD.t1195 8.10567
R306 AVDD.n1297 AVDD.t1129 8.10567
R307 AVDD.n1296 AVDD.t1013 8.10567
R308 AVDD.n1292 AVDD.t935 8.10567
R309 AVDD.n1291 AVDD.t832 8.10567
R310 AVDD.n1247 AVDD.t1245 8.10567
R311 AVDD.n1248 AVDD.t714 8.10567
R312 AVDD.n1249 AVDD.t765 8.10567
R313 AVDD.n1250 AVDD.t1169 8.10567
R314 AVDD.n1251 AVDD.t899 8.10567
R315 AVDD.n1252 AVDD.t619 8.10567
R316 AVDD.n1253 AVDD.t184 8.10567
R317 AVDD.n1254 AVDD.t237 8.10567
R318 AVDD.n1256 AVDD.t488 8.10567
R319 AVDD.n1257 AVDD.t35 8.10567
R320 AVDD.n1258 AVDD.t627 8.10567
R321 AVDD.n1259 AVDD.t204 8.10567
R322 AVDD.n1242 AVDD.t61 8.10567
R323 AVDD.n1244 AVDD.t595 8.10567
R324 AVDD.n1245 AVDD.t486 8.10567
R325 AVDD.n1302 AVDD.t563 8.10567
R326 AVDD.n1301 AVDD.t775 8.10567
R327 AVDD.n59 AVDD.t818 8.10567
R328 AVDD.n1946 AVDD.t868 8.10567
R329 AVDD.n61 AVDD.t1247 8.10567
R330 AVDD.n1941 AVDD.t995 8.10567
R331 AVDD.n62 AVDD.t731 8.10567
R332 AVDD.n1936 AVDD.t304 8.10567
R333 AVDD.n63 AVDD.t342 8.10567
R334 AVDD.n64 AVDD.t585 8.10567
R335 AVDD.n1928 AVDD.t144 8.10567
R336 AVDD.n65 AVDD.t737 8.10567
R337 AVDD.n66 AVDD.t310 8.10567
R338 AVDD.n2165 AVDD.t1111 8.10567
R339 AVDD.n30 AVDD.t852 8.10567
R340 AVDD.n2170 AVDD.t1241 8.10567
R341 AVDD.n27 AVDD.t987 8.10567
R342 AVDD.n26 AVDD.t1023 8.10567
R343 AVDD.n2177 AVDD.t609 8.10567
R344 AVDD.n1386 AVDD.t330 8.10567
R345 AVDD.n1390 AVDD.t151 8.10567
R346 AVDD.n1383 AVDD.t134 8.10567
R347 AVDD.n1395 AVDD.t548 8.10567
R348 AVDD.n1380 AVDD.t1055 8.10567
R349 AVDD.n2165 AVDD.t465 8.10567
R350 AVDD.n30 AVDD.t187 8.10567
R351 AVDD.n2170 AVDD.t617 8.10567
R352 AVDD.n27 AVDD.t340 8.10567
R353 AVDD.n26 AVDD.t375 8.10567
R354 AVDD.n2177 AVDD.t1227 8.10567
R355 AVDD.n1386 AVDD.t963 8.10567
R356 AVDD.n1390 AVDD.t812 8.10567
R357 AVDD.n1383 AVDD.t799 8.10567
R358 AVDD.n1395 AVDD.t1173 8.10567
R359 AVDD.n1380 AVDD.t411 8.10567
R360 AVDD.n501 AVDD.t735 8.10567
R361 AVDD.n502 AVDD.t1163 8.10567
R362 AVDD.n503 AVDD.t278 8.10567
R363 AVDD.n504 AVDD.t698 8.10567
R364 AVDD.n505 AVDD.t969 8.10567
R365 AVDD.n506 AVDD.t1233 8.10567
R366 AVDD.n507 AVDD.t380 8.10567
R367 AVDD.n509 AVDD.t346 8.10567
R368 AVDD.n510 AVDD.t623 8.10567
R369 AVDD.n511 AVDD.t939 8.10567
R370 AVDD.n512 AVDD.t1199 8.10567
R371 AVDD.n513 AVDD.t149 8.10567
R372 AVDD.n501 AVDD.t1139 8.10567
R373 AVDD.n502 AVDD.t290 8.10567
R374 AVDD.n503 AVDD.t674 8.10567
R375 AVDD.n504 AVDD.t1077 8.10567
R376 AVDD.n505 AVDD.t58 8.10567
R377 AVDD.n506 AVDD.t363 8.10567
R378 AVDD.n507 AVDD.t803 8.10567
R379 AVDD.n509 AVDD.t757 8.10567
R380 AVDD.n510 AVDD.t1021 8.10567
R381 AVDD.n511 AVDD.t18 8.10567
R382 AVDD.n512 AVDD.t332 8.10567
R383 AVDD.n513 AVDD.t569 8.10567
R384 AVDD.n463 AVDD.t557 8.10567
R385 AVDD.n461 AVDD.t117 8.10567
R386 AVDD.n468 AVDD.t398 8.10567
R387 AVDD.n458 AVDD.t838 8.10567
R388 AVDD.n457 AVDD.t795 8.10567
R389 AVDD.n475 AVDD.t1051 8.10567
R390 AVDD.n454 AVDD.t199 8.10567
R391 AVDD.n481 AVDD.t225 8.10567
R392 AVDD.n452 AVDD.t504 8.10567
R393 AVDD.n486 AVDD.t1029 8.10567
R394 AVDD.n449 AVDD.t1279 8.10567
R395 AVDD.n463 AVDD.t949 8.10567
R396 AVDD.n461 AVDD.t522 8.10567
R397 AVDD.n468 AVDD.t814 8.10567
R398 AVDD.n458 AVDD.t1217 8.10567
R399 AVDD.n457 AVDD.t1175 8.10567
R400 AVDD.n475 AVDD.t173 8.10567
R401 AVDD.n454 AVDD.t611 8.10567
R402 AVDD.n481 AVDD.t629 8.10567
R403 AVDD.n452 AVDD.t915 8.10567
R404 AVDD.n486 AVDD.t146 8.10567
R405 AVDD.n449 AVDD.t433 8.10567
R406 AVDD.n519 AVDD.t1255 8.10567
R407 AVDD.n518 AVDD.t99 8.10567
R408 AVDD.n602 AVDD.t66 8.10567
R409 AVDD.n601 AVDD.t202 8.10567
R410 AVDD.n599 AVDD.t979 8.10567
R411 AVDD.n612 AVDD.t1093 8.10567
R412 AVDD.n611 AVDD.t997 8.10567
R413 AVDD.n515 AVDD.t1003 8.10567
R414 AVDD.n516 AVDD.t635 8.10567
R415 AVDD.n1466 AVDD.t453 8.10567
R416 AVDD.n670 AVDD.t1039 8.10567
R417 AVDD.n1471 AVDD.t1109 8.10567
R418 AVDD.n667 AVDD.t761 8.10567
R419 AVDD.n124 AVDD.t154 8.10567
R420 AVDD.n1478 AVDD.t230 8.10567
R421 AVDD.n664 AVDD.t1145 8.10567
R422 AVDD.n125 AVDD.t461 8.10567
R423 AVDD.n126 AVDD.t534 8.10567
R424 AVDD.n127 AVDD.t163 8.10567
R425 AVDD.n128 AVDD.t243 8.10567
R426 AVDD.n129 AVDD.t967 8.10567
R427 AVDD.n134 AVDD.t407 8.10567
R428 AVDD.n135 AVDD.t1147 8.10567
R429 AVDD.n136 AVDD.t785 8.10567
R430 AVDD.n137 AVDD.t856 8.10567
R431 AVDD.n138 AVDD.t459 8.10567
R432 AVDD.n139 AVDD.t858 8.10567
R433 AVDD.n140 AVDD.t907 8.10567
R434 AVDD.n141 AVDD.t530 8.10567
R435 AVDD.n143 AVDD.t1223 8.10567
R436 AVDD.n144 AVDD.t1269 8.10567
R437 AVDD.n145 AVDD.t767 8.10567
R438 AVDD.n146 AVDD.t820 8.10567
R439 AVDD.n147 AVDD.t591 8.10567
R440 AVDD.n1466 AVDD.t463 8.10567
R441 AVDD.n670 AVDD.t1047 8.10567
R442 AVDD.n1471 AVDD.t1117 8.10567
R443 AVDD.n667 AVDD.t769 8.10567
R444 AVDD.n124 AVDD.t159 8.10567
R445 AVDD.n1478 AVDD.t235 8.10567
R446 AVDD.n664 AVDD.t1151 8.10567
R447 AVDD.n125 AVDD.t473 8.10567
R448 AVDD.n126 AVDD.t540 8.10567
R449 AVDD.n127 AVDD.t171 8.10567
R450 AVDD.n128 AVDD.t249 8.10567
R451 AVDD.n129 AVDD.t975 8.10567
R452 AVDD.n134 AVDD.t409 8.10567
R453 AVDD.n135 AVDD.t1155 8.10567
R454 AVDD.n136 AVDD.t787 8.10567
R455 AVDD.n137 AVDD.t864 8.10567
R456 AVDD.n138 AVDD.t467 8.10567
R457 AVDD.n139 AVDD.t860 8.10567
R458 AVDD.n140 AVDD.t913 8.10567
R459 AVDD.n141 AVDD.t538 8.10567
R460 AVDD.n143 AVDD.t1229 8.10567
R461 AVDD.n144 AVDD.t1273 8.10567
R462 AVDD.n145 AVDD.t771 8.10567
R463 AVDD.n146 AVDD.t828 8.10567
R464 AVDD.n147 AVDD.t597 8.10567
R465 AVDD.n490 AVDD.t197 8.10567
R466 AVDD.n491 AVDD.t55 8.10567
R467 AVDD.n496 AVDD.t74 8.10567
R468 AVDD.n497 AVDD.t546 8.10567
R469 AVDD.n499 AVDD.t603 8.10567
R470 AVDD.n490 AVDD.t929 8.10567
R471 AVDD.n491 AVDD.t824 8.10567
R472 AVDD.n496 AVDD.t842 8.10567
R473 AVDD.n497 AVDD.t830 8.10567
R474 AVDD.n499 AVDD.t161 8.10567
R475 AVDD.n556 AVDD.t1001 8.10567
R476 AVDD.n558 AVDD.t419 8.10567
R477 AVDD.n559 AVDD.t544 8.10567
R478 AVDD.n564 AVDD.t528 8.10567
R479 AVDD.n565 AVDD.t633 8.10567
R480 AVDD.n567 AVDD.t125 8.10567
R481 AVDD.n556 AVDD.t581 8.10567
R482 AVDD.n558 AVDD.t1257 8.10567
R483 AVDD.n559 AVDD.t107 8.10567
R484 AVDD.n564 AVDD.t78 8.10567
R485 AVDD.n565 AVDD.t213 8.10567
R486 AVDD.n567 AVDD.t989 8.10567
R487 AVDD.n571 AVDD.t274 8.10567
R488 AVDD.n415 AVDD.t688 8.10567
R489 AVDD.n576 AVDD.t1061 8.10567
R490 AVDD.n414 AVDD.t217 8.10567
R491 AVDD.n413 AVDD.t490 8.10567
R492 AVDD.n583 AVDD.t791 8.10567
R493 AVDD.n412 AVDD.t1189 8.10567
R494 AVDD.n589 AVDD.t1159 8.10567
R495 AVDD.n411 AVDD.t132 8.10567
R496 AVDD.n594 AVDD.t445 8.10567
R497 AVDD.n410 AVDD.t749 8.10567
R498 AVDD.n422 AVDD.t50 8.10567
R499 AVDD.n421 AVDD.t943 8.10567
R500 AVDD.n427 AVDD.t1201 8.10567
R501 AVDD.n420 AVDD.t359 8.10567
R502 AVDD.n419 AVDD.t316 8.10567
R503 AVDD.n434 AVDD.t589 8.10567
R504 AVDD.n418 AVDD.t1011 8.10567
R505 AVDD.n440 AVDD.t1027 8.10567
R506 AVDD.n417 AVDD.t1277 8.10567
R507 AVDD.n445 AVDD.t579 8.10567
R508 AVDD.n416 AVDD.t872 8.10567
R509 AVDD.n1484 AVDD.t209 8.10567
R510 AVDD.n1486 AVDD.t729 8.10567
R511 AVDD.n1487 AVDD.t607 8.10567
R512 AVDD.n1492 AVDD.t684 8.10567
R513 AVDD.n1491 AVDD.t893 8.10567
R514 AVDD.n1489 AVDD.t94 8.10567
R515 AVDD.n1484 AVDD.t1049 8.10567
R516 AVDD.n1486 AVDD.t300 8.10567
R517 AVDD.n1487 AVDD.t165 8.10567
R518 AVDD.n1492 AVDD.t270 8.10567
R519 AVDD.n1491 AVDD.t439 8.10567
R520 AVDD.n1489 AVDD.t957 8.10567
R521 AVDD.n1503 AVDD.t753 8.10567
R522 AVDD.n1501 AVDD.t1237 8.10567
R523 AVDD.n1500 AVDD.t1143 8.10567
R524 AVDD.n130 AVDD.t498 8.10567
R525 AVDD.n131 AVDD.t389 8.10567
R526 AVDD.n1503 AVDD.t318 8.10567
R527 AVDD.n1501 AVDD.t836 8.10567
R528 AVDD.n1500 AVDD.t721 8.10567
R529 AVDD.n130 AVDD.t1219 8.10567
R530 AVDD.n131 AVDD.t1115 8.10567
R531 AVDD.n1507 AVDD.t240 8.10567
R532 AVDD.n107 AVDD.t660 8.10567
R533 AVDD.n1512 AVDD.t1033 8.10567
R534 AVDD.n104 AVDD.t191 8.10567
R535 AVDD.n103 AVDD.t455 8.10567
R536 AVDD.n1519 AVDD.t763 8.10567
R537 AVDD.n381 AVDD.t1171 8.10567
R538 AVDD.n385 AVDD.t1127 8.10567
R539 AVDD.n378 AVDD.t120 8.10567
R540 AVDD.n390 AVDD.t423 8.10567
R541 AVDD.n375 AVDD.t727 8.10567
R542 AVDD.n395 AVDD.t951 8.10567
R543 AVDD.n1507 AVDD.t885 8.10567
R544 AVDD.n107 AVDD.t1267 8.10567
R545 AVDD.n1512 AVDD.t403 8.10567
R546 AVDD.n104 AVDD.t846 8.10567
R547 AVDD.n103 AVDD.t1091 8.10567
R548 AVDD.n1519 AVDD.t86 8.10567
R549 AVDD.n381 AVDD.t524 8.10567
R550 AVDD.n385 AVDD.t482 8.10567
R551 AVDD.n378 AVDD.t777 8.10567
R552 AVDD.n390 AVDD.t1057 8.10567
R553 AVDD.n375 AVDD.t43 8.10567
R554 AVDD.n395 AVDD.t308 8.10567
R555 AVDD.n398 AVDD.t822 8.10567
R556 AVDD.n399 AVDD.t710 8.10567
R557 AVDD.n404 AVDD.t123 8.10567
R558 AVDD.n405 AVDD.t1271 8.10567
R559 AVDD.n363 AVDD.t1037 8.10567
R560 AVDD.n365 AVDD.t296 8.10567
R561 AVDD.n366 AVDD.t157 8.10567
R562 AVDD.n371 AVDD.t259 8.10567
R563 AVDD.n372 AVDD.t427 8.10567
R564 AVDD.n86 AVDD.t344 8.10567
R565 AVDD.n1535 AVDD.t779 8.10567
R566 AVDD.n88 AVDD.t1161 8.10567
R567 AVDD.n1530 AVDD.t306 8.10567
R568 AVDD.n89 AVDD.t575 8.10567
R569 AVDD.n1525 AVDD.t870 8.10567
R570 AVDD.n349 AVDD.t1253 8.10567
R571 AVDD.n353 AVDD.t1213 8.10567
R572 AVDD.n348 AVDD.t223 8.10567
R573 AVDD.n358 AVDD.t536 8.10567
R574 AVDD.n150 AVDD.t826 8.10567
R575 AVDD.n1399 AVDD.t21 8.10567
R576 AVDD.n1400 AVDD.t917 8.10567
R577 AVDD.n1401 AVDD.t1181 8.10567
R578 AVDD.n1402 AVDD.t337 8.10567
R579 AVDD.n1403 AVDD.t298 8.10567
R580 AVDD.n1404 AVDD.t567 8.10567
R581 AVDD.n1405 AVDD.t993 8.10567
R582 AVDD.n1406 AVDD.t1009 8.10567
R583 AVDD.n1407 AVDD.t1265 8.10567
R584 AVDD.n1408 AVDD.t559 8.10567
R585 AVDD.n1409 AVDD.t844 8.10567
R586 AVDD.n1399 AVDD.t692 8.10567
R587 AVDD.n1400 AVDD.t276 8.10567
R588 AVDD.n1401 AVDD.t552 8.10567
R589 AVDD.n1402 AVDD.t973 8.10567
R590 AVDD.n1403 AVDD.t927 8.10567
R591 AVDD.n1404 AVDD.t1193 8.10567
R592 AVDD.n1405 AVDD.t351 8.10567
R593 AVDD.n1406 AVDD.t368 8.10567
R594 AVDD.n1407 AVDD.t648 8.10567
R595 AVDD.n1408 AVDD.t1179 8.10567
R596 AVDD.n1409 AVDD.t176 8.10567
R597 AVDD.n1029 AVDD.t1079 8.10567
R598 AVDD.n1001 AVDD.t658 8.10567
R599 AVDD.n957 AVDD.t783 8.10567
R600 AVDD.n990 AVDD.t189 8.10567
R601 AVDD.n1203 AVDD.t945 8.10567
R602 AVDD.n1202 AVDD.t129 8.10567
R603 AVDD.n717 AVDD.t678 8.10567
R604 AVDD.n1223 AVDD.t1185 8.10567
R605 AVDD.n769 AVDD.t921 8.10567
R606 AVDD.n773 AVDD.t640 8.10567
R607 AVDD.n763 AVDD.t215 8.10567
R608 AVDD.n758 AVDD.t272 8.10567
R609 AVDD.n946 AVDD.t510 8.10567
R610 AVDD.n755 AVDD.t64 8.10567
R611 AVDD.n783 AVDD.t656 8.10567
R612 AVDD.n782 AVDD.t228 8.10567
R613 AVDD.n786 AVDD.t1249 8.10567
R614 AVDD.n904 AVDD.t76 8.10567
R615 AVDD.n920 AVDD.t1153 8.10567
R616 AVDD.n917 AVDD.t879 8.10567
R617 AVDD.n1225 AVDD.t654 8.10567
R618 AVDD.n767 AVDD.t1203 8.10567
R619 AVDD.n774 AVDD.t743 8.10567
R620 AVDD.n759 AVDD.t365 8.10567
R621 AVDD.n760 AVDD.t1251 8.10567
R622 AVDD.n947 AVDD.t1043 8.10567
R623 AVDD.n754 AVDD.t1121 8.10567
R624 AVDD.n784 AVDD.t26 8.10567
R625 AVDD.n785 AVDD.t686 8.10567
R626 AVDD.n933 AVDD.t901 8.10567
R627 AVDD.n905 AVDD.t961 8.10567
R628 AVDD.n926 AVDD.t475 8.10567
R629 AVDD.n921 AVDD.t615 8.10567
R630 AVDD.n712 AVDD.t739 8.10567
R631 AVDD.n1230 AVDD.t789 8.10567
R632 AVDD.n803 AVDD.t312 8.10567
R633 AVDD.n802 AVDD.t413 8.10567
R634 AVDD.n1238 AVDD.t405 8.10567
R635 AVDD.n1237 AVDD.t516 8.10567
R636 AVDD.n1235 AVDD.t1261 8.10567
R637 AVDD.n915 AVDD.t1259 8.10567
R638 AVDD.n907 AVDD.t1005 8.10567
R639 AVDD.n908 AVDD.t1041 8.10567
R640 AVDD.n19 AVDD.t631 8.10567
R641 AVDD.n18 AVDD.t355 8.10567
R642 AVDD.n2187 AVDD.t182 8.10567
R643 AVDD.n17 AVDD.t169 8.10567
R644 AVDD.n2192 AVDD.t571 8.10567
R645 AVDD.n16 AVDD.t1073 8.10567
R646 AVDD.n880 AVDD.t565 8.10567
R647 AVDD.n881 AVDD.t437 8.10567
R648 AVDD.n886 AVDD.t449 8.10567
R649 AVDD.n887 AVDD.t1017 8.10567
R650 AVDD.n889 AVDD.t447 8.10567
R651 AVDD.n880 AVDD.t142 8.10567
R652 AVDD.n881 AVDD.t15 8.10567
R653 AVDD.n886 AVDD.t41 8.10567
R654 AVDD.n887 AVDD.t700 8.10567
R655 AVDD.n889 AVDD.t573 8.10567
R656 AVDD.n893 AVDD.t877 8.10567
R657 AVDD.n895 AVDD.t302 8.10567
R658 AVDD.n896 AVDD.t401 8.10567
R659 AVDD.n900 AVDD.t385 8.10567
R660 AVDD.n901 AVDD.t496 8.10567
R661 AVDD.n893 AVDD.t977 8.10567
R662 AVDD.n895 AVDD.t396 8.10567
R663 AVDD.n896 AVDD.t512 8.10567
R664 AVDD.n900 AVDD.t492 8.10567
R665 AVDD.n901 AVDD.t613 8.10567
R666 AVDD.n839 AVDD.t334 8.10567
R667 AVDD.n840 AVDD.t29 8.10567
R668 AVDD.n841 AVDD.t469 8.10567
R669 AVDD.n842 AVDD.t194 8.10567
R670 AVDD.n843 AVDD.t251 8.10567
R671 AVDD.n844 AVDD.t1085 8.10567
R672 AVDD.n845 AVDD.t834 8.10567
R673 AVDD.n847 AVDD.t662 8.10567
R674 AVDD.n848 AVDD.t644 8.10567
R675 AVDD.n849 AVDD.t1025 8.10567
R676 AVDD.n850 AVDD.t293 8.10567
R677 AVDD.n839 AVDD.t745 8.10567
R678 AVDD.n840 AVDD.t443 8.10567
R679 AVDD.n841 AVDD.t891 8.10567
R680 AVDD.n842 AVDD.t601 8.10567
R681 AVDD.n843 AVDD.t646 8.10567
R682 AVDD.n844 AVDD.t219 8.10567
R683 AVDD.n845 AVDD.t1211 8.10567
R684 AVDD.n847 AVDD.t1053 8.10567
R685 AVDD.n848 AVDD.t1031 8.10567
R686 AVDD.n849 AVDD.t139 8.10567
R687 AVDD.n850 AVDD.t682 8.10567
R688 AVDD.n801 AVDD.t477 8.10567
R689 AVDD.n812 AVDD.t1197 8.10567
R690 AVDD.n799 AVDD.t1231 8.10567
R691 AVDD.n817 AVDD.t377 8.10567
R692 AVDD.n796 AVDD.t91 8.10567
R693 AVDD.n795 AVDD.t1101 8.10567
R694 AVDD.n824 AVDD.t696 8.10567
R695 AVDD.n792 AVDD.t733 8.10567
R696 AVDD.n830 AVDD.t985 8.10567
R697 AVDD.n790 AVDD.t561 8.10567
R698 AVDD.n835 AVDD.t1123 8.10567
R699 AVDD.n787 AVDD.t708 8.10567
R700 AVDD.n801 AVDD.t895 8.10567
R701 AVDD.n812 AVDD.t325 8.10567
R702 AVDD.n799 AVDD.t361 8.10567
R703 AVDD.n817 AVDD.t801 8.10567
R704 AVDD.n796 AVDD.t506 8.10567
R705 AVDD.n795 AVDD.t232 8.10567
R706 AVDD.n824 AVDD.t1071 8.10567
R707 AVDD.n792 AVDD.t1137 8.10567
R708 AVDD.n830 AVDD.t81 8.10567
R709 AVDD.n790 AVDD.t955 8.10567
R710 AVDD.n835 AVDD.t254 8.10567
R711 AVDD.n787 AVDD.t1087 8.10567
R712 AVDD.n741 AVDD.t983 8.10567
R713 AVDD.n742 AVDD.t179 8.10567
R714 AVDD.n1180 AVDD.t723 8.10567
R715 AVDD.n1007 AVDD.t1141 8.10567
R716 AVDD.n1009 AVDD.t706 8.10567
R717 AVDD.n1008 AVDD.t816 8.10567
R718 AVDD.n1097 AVDD.t245 8.10567
R719 AVDD.n983 AVDD.t809 8.10567
R720 AVDD.n1092 AVDD.t322 8.10567
R721 AVDD.n984 AVDD.t1221 8.10567
R722 AVDD.n1087 AVDD.t874 8.10567
R723 AVDD.n985 AVDD.t637 8.10567
R724 AVDD.n1082 AVDD.t716 8.10567
R725 AVDD.n986 AVDD.t925 8.10567
R726 AVDD.n987 AVDD.t281 8.10567
R727 AVDD.n1074 AVDD.t479 8.10567
R728 AVDD.n988 AVDD.t554 8.10567
R729 AVDD.n1069 AVDD.t38 8.10567
R730 AVDD.n1247 AVDD.t621 8.10567
R731 AVDD.n1248 AVDD.t32 8.10567
R732 AVDD.n1249 AVDD.t84 8.10567
R733 AVDD.n1250 AVDD.t518 8.10567
R734 AVDD.n1251 AVDD.t257 8.10567
R735 AVDD.n1252 AVDD.t1239 8.10567
R736 AVDD.n1253 AVDD.t840 8.10567
R737 AVDD.n1254 AVDD.t883 8.10567
R738 AVDD.n1256 AVDD.t1113 8.10567
R739 AVDD.n1257 AVDD.t704 8.10567
R740 AVDD.n1258 AVDD.t1243 8.10567
R741 AVDD.n1259 AVDD.t850 8.10567
R742 AVDD.n999 AVDD.t327 6.64567
R743 AVDD.n1036 AVDD.t393 6.64567
R744 AVDD.n997 AVDD.t1183 6.64567
R745 AVDD.n996 AVDD.t991 6.64567
R746 AVDD.n1043 AVDD.t1275 6.64567
R747 AVDD.n1045 AVDD.t919 6.64567
R748 AVDD.n1046 AVDD.t542 6.64567
R749 AVDD.n1046 AVDD.t887 6.64567
R750 AVDD.n1052 AVDD.t807 6.64567
R751 AVDD.n1052 AVDD.t1131 6.64567
R752 AVDD.n1053 AVDD.t435 6.64567
R753 AVDD.n1053 AVDD.t797 6.64567
R754 AVDD.n1055 AVDD.t1 6.64567
R755 AVDD.n1055 AVDD.t372 6.64567
R756 AVDD.n993 AVDD.t666 6.64567
R757 AVDD.n1062 AVDD.t741 6.64567
R758 AVDD.n1058 AVDD.t263 6.64567
R759 AVDD.n1030 AVDD.t12 6.64567
R760 AVDD.n1004 AVDD.t931 6.64567
R761 AVDD.n1002 AVDD.t897 6.64567
R762 AVDD.n1118 AVDD.t1149 6.64567
R763 AVDD.n958 AVDD.t805 6.64567
R764 AVDD.n991 AVDD.t387 6.64567
R765 AVDD.n1920 AVDD.t1900 6.58663
R766 AVDD.n1852 AVDD.t1541 6.58663
R767 AVDD.n154 AVDD.t1813 6.58663
R768 AVDD.n262 AVDD.t1397 6.58663
R769 AVDD.n2115 AVDD.n2109 6.50088
R770 AVDD.n2048 AVDD.n2047 6.50088
R771 AVDD.n1706 AVDD.n1705 6.50088
R772 AVDD.n1647 AVDD.n1641 6.50088
R773 AVDD.n1857 AVDD.n1856 6.45575
R774 AVDD.n1790 AVDD.n1782 6.45575
R775 AVDD.n289 AVDD.n280 6.45575
R776 AVDD.n232 AVDD.n223 6.45575
R777 AVDD.n1921 AVDD.n1917 5.95439
R778 AVDD.n1853 AVDD.n1849 5.95439
R779 AVDD.n342 AVDD.n341 5.95439
R780 AVDD.n264 AVDD.n263 5.95439
R781 AVDD.n1917 AVDD.t1651 5.31528
R782 AVDD.n1849 AVDD.t1584 5.31528
R783 AVDD.n342 AVDD.t1764 5.31528
R784 AVDD.n264 AVDD.t1357 5.31528
R785 AVDD.n1057 AVDD.n995 5.19255
R786 AVDD.n1215 AVDD.t1529 5.12594
R787 AVDD.n1496 AVDD.n114 5.12014
R788 AVDD.n2154 AVDD.n37 5.12014
R789 AVDD.n1018 AVDD.t1293 5.09041
R790 AVDD.t329 AVDD.n1033 5.0505
R791 AVDD.n1039 AVDD.t1184 5.0505
R792 AVDD.t992 AVDD.n1040 5.0505
R793 AVDD.n1041 AVDD.t992 5.0505
R794 AVDD.t265 AVDD.n1059 5.0505
R795 AVDD.n1065 AVDD.t667 5.0505
R796 AVDD.n1779 AVDD.n1778 4.96877
R797 AVDD.n1771 AVDD.n1770 4.96877
R798 AVDD.n229 AVDD.n228 4.96877
R799 AVDD.n286 AVDD.n285 4.96877
R800 AVDD.n51 AVDD.n48 4.92758
R801 AVDD.n2054 AVDD.n2051 4.92758
R802 AVDD.n78 AVDD.n75 4.92758
R803 AVDD.n1655 AVDD.n1652 4.92758
R804 AVDD.n1962 AVDD.n1961 4.78594
R805 AVDD.n1985 AVDD.n1984 4.78594
R806 AVDD.n1547 AVDD.n1546 4.78594
R807 AVDD.n1594 AVDD.n1593 4.78594
R808 AVDD.n1780 AVDD.n1779 4.61712
R809 AVDD.n1794 AVDD.n1793 4.61712
R810 AVDD.n1772 AVDD.n1771 4.61712
R811 AVDD.n1861 AVDD.n1860 4.61712
R812 AVDD.n230 AVDD.n229 4.61712
R813 AVDD.n217 AVDD.n216 4.61712
R814 AVDD.n287 AVDD.n286 4.61712
R815 AVDD.n274 AVDD.n273 4.61712
R816 AVDD.n2099 AVDD.n2095 4.61078
R817 AVDD.n2093 AVDD.n2089 4.61078
R818 AVDD.n2087 AVDD.n2083 4.61078
R819 AVDD.n2081 AVDD.n2077 4.61078
R820 AVDD.n1978 AVDD.n1974 4.61078
R821 AVDD.n1972 AVDD.n1968 4.61078
R822 AVDD.n1966 AVDD.n1962 4.61078
R823 AVDD.n2037 AVDD.n2033 4.61078
R824 AVDD.n2031 AVDD.n2027 4.61078
R825 AVDD.n2025 AVDD.n2021 4.61078
R826 AVDD.n2019 AVDD.n2015 4.61078
R827 AVDD.n2001 AVDD.n1997 4.61078
R828 AVDD.n1995 AVDD.n1991 4.61078
R829 AVDD.n1989 AVDD.n1985 4.61078
R830 AVDD.n1792 AVDD.n1791 4.61078
R831 AVDD.n1859 AVDD.n1858 4.61078
R832 AVDD.n1679 AVDD.n1678 4.61078
R833 AVDD.n1682 AVDD.n1681 4.61078
R834 AVDD.n1685 AVDD.n1684 4.61078
R835 AVDD.n1688 AVDD.n1687 4.61078
R836 AVDD.n1563 AVDD.n1559 4.61078
R837 AVDD.n1557 AVDD.n1553 4.61078
R838 AVDD.n1551 AVDD.n1547 4.61078
R839 AVDD.n1629 AVDD.n1628 4.61078
R840 AVDD.n1632 AVDD.n1631 4.61078
R841 AVDD.n1635 AVDD.n1634 4.61078
R842 AVDD.n1638 AVDD.n1637 4.61078
R843 AVDD.n1610 AVDD.n1606 4.61078
R844 AVDD.n1604 AVDD.n1600 4.61078
R845 AVDD.n1598 AVDD.n1594 4.61078
R846 AVDD.n222 AVDD.n218 4.61078
R847 AVDD.n279 AVDD.n275 4.61078
R848 AVDD.n1176 AVDD.n1170 4.61078
R849 AVDD.n1168 AVDD.n1162 4.61078
R850 AVDD.n1160 AVDD.n1154 4.61078
R851 AVDD.n1152 AVDD.n1148 4.61078
R852 AVDD.n1146 AVDD.n1140 4.61078
R853 AVDD.n1138 AVDD.n1132 4.61078
R854 AVDD.n1101 AVDD.n1100 4.61078
R855 AVDD.n1104 AVDD.n1103 4.61078
R856 AVDD.n1107 AVDD.n1106 4.61078
R857 AVDD.n1110 AVDD.n1109 4.61078
R858 AVDD.n1113 AVDD.n1112 4.61078
R859 AVDD.n1116 AVDD.n1115 4.61078
R860 AVDD.n1184 AVDD.n1183 4.60951
R861 AVDD.n1183 AVDD.n1182 4.60951
R862 AVDD.n1187 AVDD.n1186 4.60951
R863 AVDD.n1186 AVDD.n1185 4.60951
R864 AVDD.n1190 AVDD.n1189 4.60951
R865 AVDD.n1189 AVDD.n1188 4.60951
R866 AVDD.n1193 AVDD.n1192 4.60951
R867 AVDD.n1192 AVDD.n1191 4.60951
R868 AVDD.n1196 AVDD.n1195 4.60951
R869 AVDD.n1195 AVDD.n1194 4.60951
R870 AVDD.n1199 AVDD.n1198 4.60951
R871 AVDD.n1198 AVDD.n1197 4.60951
R872 AVDD.n2100 AVDD.n2099 4.60825
R873 AVDD.n2094 AVDD.n2093 4.60825
R874 AVDD.n2088 AVDD.n2087 4.60825
R875 AVDD.n2082 AVDD.n2081 4.60825
R876 AVDD.n1979 AVDD.n1978 4.60825
R877 AVDD.n1973 AVDD.n1972 4.60825
R878 AVDD.n1967 AVDD.n1966 4.60825
R879 AVDD.n2038 AVDD.n2037 4.60825
R880 AVDD.n2032 AVDD.n2031 4.60825
R881 AVDD.n2026 AVDD.n2025 4.60825
R882 AVDD.n2020 AVDD.n2019 4.60825
R883 AVDD.n2002 AVDD.n2001 4.60825
R884 AVDD.n1996 AVDD.n1995 4.60825
R885 AVDD.n1990 AVDD.n1989 4.60825
R886 AVDD.n1791 AVDD.n1790 4.60825
R887 AVDD.n1858 AVDD.n1857 4.60825
R888 AVDD.n1678 AVDD.n1677 4.60825
R889 AVDD.n1681 AVDD.n1680 4.60825
R890 AVDD.n1684 AVDD.n1683 4.60825
R891 AVDD.n1687 AVDD.n1686 4.60825
R892 AVDD.n1564 AVDD.n1563 4.60825
R893 AVDD.n1558 AVDD.n1557 4.60825
R894 AVDD.n1552 AVDD.n1551 4.60825
R895 AVDD.n1628 AVDD.n1581 4.60825
R896 AVDD.n1631 AVDD.n1630 4.60825
R897 AVDD.n1634 AVDD.n1633 4.60825
R898 AVDD.n1637 AVDD.n1636 4.60825
R899 AVDD.n1611 AVDD.n1610 4.60825
R900 AVDD.n1605 AVDD.n1604 4.60825
R901 AVDD.n1599 AVDD.n1598 4.60825
R902 AVDD.n223 AVDD.n222 4.60825
R903 AVDD.n280 AVDD.n279 4.60825
R904 AVDD.n1177 AVDD.n1176 4.60825
R905 AVDD.n1169 AVDD.n1168 4.60825
R906 AVDD.n1161 AVDD.n1160 4.60825
R907 AVDD.n1153 AVDD.n1152 4.60825
R908 AVDD.n1147 AVDD.n1146 4.60825
R909 AVDD.n1139 AVDD.n1138 4.60825
R910 AVDD.n1100 AVDD.n1099 4.60825
R911 AVDD.n1103 AVDD.n1102 4.60825
R912 AVDD.n1106 AVDD.n1105 4.60825
R913 AVDD.n1109 AVDD.n1108 4.60825
R914 AVDD.n1112 AVDD.n1111 4.60825
R915 AVDD.n1115 AVDD.n1114 4.60825
R916 AVDD.n1781 AVDD.n1780 4.60191
R917 AVDD.n1795 AVDD.n1794 4.60191
R918 AVDD.n1773 AVDD.n1772 4.60191
R919 AVDD.n1862 AVDD.n1861 4.60191
R920 AVDD.n231 AVDD.n230 4.60191
R921 AVDD.n216 AVDD.n188 4.60191
R922 AVDD.n288 AVDD.n287 4.60191
R923 AVDD.n273 AVDD.n270 4.60191
R924 AVDD.n1916 AVDD.n1913 4.50663
R925 AVDD.n1848 AVDD.n1758 4.50663
R926 AVDD.n346 AVDD.n345 4.50663
R927 AVDD.n268 AVDD.n267 4.50663
R928 AVDD.n1965 AVDD.n1959 4.5005
R929 AVDD.n1971 AVDD.n1958 4.5005
R930 AVDD.n1977 AVDD.n1957 4.5005
R931 AVDD.n2080 AVDD.n1956 4.5005
R932 AVDD.n2086 AVDD.n1955 4.5005
R933 AVDD.n2092 AVDD.n1954 4.5005
R934 AVDD.n2098 AVDD.n1953 4.5005
R935 AVDD.n1988 AVDD.n1982 4.5005
R936 AVDD.n1994 AVDD.n1981 4.5005
R937 AVDD.n2000 AVDD.n1980 4.5005
R938 AVDD.n2018 AVDD.n2014 4.5005
R939 AVDD.n2024 AVDD.n2013 4.5005
R940 AVDD.n2030 AVDD.n2012 4.5005
R941 AVDD.n2036 AVDD.n2011 4.5005
R942 AVDD.n1761 AVDD.n1759 4.5005
R943 AVDD.n1765 AVDD.n1762 4.5005
R944 AVDD.n1768 AVDD.n1766 4.5005
R945 AVDD.n1785 AVDD.n1783 4.5005
R946 AVDD.n1789 AVDD.n1786 4.5005
R947 AVDD.n1776 AVDD.n1774 4.5005
R948 AVDD.n1550 AVDD.n1544 4.5005
R949 AVDD.n1556 AVDD.n1543 4.5005
R950 AVDD.n1562 AVDD.n1542 4.5005
R951 AVDD.n1568 AVDD.n1565 4.5005
R952 AVDD.n1572 AVDD.n1569 4.5005
R953 AVDD.n1576 AVDD.n1573 4.5005
R954 AVDD.n1580 AVDD.n1577 4.5005
R955 AVDD.n1597 AVDD.n1591 4.5005
R956 AVDD.n1603 AVDD.n1590 4.5005
R957 AVDD.n1609 AVDD.n1589 4.5005
R958 AVDD.n1615 AVDD.n1612 4.5005
R959 AVDD.n1619 AVDD.n1616 4.5005
R960 AVDD.n1623 AVDD.n1620 4.5005
R961 AVDD.n1627 AVDD.n1624 4.5005
R962 AVDD.n272 AVDD.n187 4.5005
R963 AVDD.n278 AVDD.n186 4.5005
R964 AVDD.n283 AVDD.n281 4.5005
R965 AVDD.n215 AVDD.n213 4.5005
R966 AVDD.n221 AVDD.n212 4.5005
R967 AVDD.n226 AVDD.n224 4.5005
R968 AVDD.n721 AVDD.n718 4.5005
R969 AVDD.n725 AVDD.n722 4.5005
R970 AVDD.n728 AVDD.n726 4.5005
R971 AVDD.n732 AVDD.n729 4.5005
R972 AVDD.n736 AVDD.n733 4.5005
R973 AVDD.n740 AVDD.n737 4.5005
R974 AVDD.n1135 AVDD.n750 4.5005
R975 AVDD.n1143 AVDD.n749 4.5005
R976 AVDD.n1150 AVDD.n748 4.5005
R977 AVDD.n1157 AVDD.n747 4.5005
R978 AVDD.n1165 AVDD.n746 4.5005
R979 AVDD.n1173 AVDD.n745 4.5005
R980 AVDD.n962 AVDD.n959 4.5005
R981 AVDD.n966 AVDD.n963 4.5005
R982 AVDD.n969 AVDD.n967 4.5005
R983 AVDD.n973 AVDD.n970 4.5005
R984 AVDD.n977 AVDD.n974 4.5005
R985 AVDD.n981 AVDD.n978 4.5005
R986 AVDD.n1796 AVDD.n1795 4.32507
R987 AVDD.n259 AVDD.n188 4.32507
R988 AVDD.n2040 AVDD.t1649 4.06712
R989 AVDD.n2009 AVDD.t1607 4.06712
R990 AVDD.n2116 AVDD.t1290 4.06712
R991 AVDD.n2107 AVDD.t1326 4.06712
R992 AVDD.n1648 AVDD.t1415 4.06712
R993 AVDD.n1587 AVDD.t1384 4.06712
R994 AVDD.n1698 AVDD.t1836 4.06712
R995 AVDD.n1696 AVDD.t1791 4.06712
R996 AVDD.n2118 AVDD.n2117 3.96014
R997 AVDD.n2041 AVDD.n2039 3.96014
R998 AVDD.n1699 AVDD.n73 3.96014
R999 AVDD.n1650 AVDD.n1649 3.96014
R1000 AVDD.n2040 AVDD.t1499 3.86107
R1001 AVDD.n2009 AVDD.t1671 3.86107
R1002 AVDD.n2116 AVDD.t1869 3.86107
R1003 AVDD.n2107 AVDD.t1317 3.86107
R1004 AVDD.n1648 AVDD.t1789 3.86107
R1005 AVDD.n1587 AVDD.t1344 3.86107
R1006 AVDD.n1698 AVDD.t1822 3.86107
R1007 AVDD.n1696 AVDD.t1776 3.86107
R1008 AVDD.n1776 AVDD.n1775 3.84568
R1009 AVDD.n1785 AVDD.n1784 3.84568
R1010 AVDD.n1768 AVDD.n1767 3.84568
R1011 AVDD.n1761 AVDD.n1760 3.84568
R1012 AVDD.n226 AVDD.n225 3.84568
R1013 AVDD.n215 AVDD.n214 3.84568
R1014 AVDD.n283 AVDD.n282 3.84568
R1015 AVDD.n272 AVDD.n271 3.84568
R1016 AVDD.n1920 AVDD.n1919 3.84528
R1017 AVDD.n1916 AVDD.n1915 3.84528
R1018 AVDD.n1852 AVDD.n1851 3.84528
R1019 AVDD.n1848 AVDD.n1847 3.84528
R1020 AVDD.n154 AVDD.n153 3.84528
R1021 AVDD.n345 AVDD.n344 3.84528
R1022 AVDD.n262 AVDD.n261 3.84528
R1023 AVDD.n267 AVDD.n266 3.84528
R1024 AVDD.n1152 AVDD.n1151 3.84449
R1025 AVDD.n54 AVDD.n51 3.79678
R1026 AVDD.n2128 AVDD.n2125 3.79678
R1027 AVDD.n2057 AVDD.n2054 3.79678
R1028 AVDD.n2069 AVDD.n2066 3.79678
R1029 AVDD.n1905 AVDD.n1899 3.79678
R1030 AVDD.n1880 AVDD.n1874 3.79678
R1031 AVDD.n1814 AVDD.n1808 3.79678
R1032 AVDD.n1837 AVDD.n1831 3.79678
R1033 AVDD.n81 AVDD.n78 3.79678
R1034 AVDD.n1718 AVDD.n1715 3.79678
R1035 AVDD.n1658 AVDD.n1655 3.79678
R1036 AVDD.n1671 AVDD.n1668 3.79678
R1037 AVDD.n308 AVDD.n302 3.79678
R1038 AVDD.n331 AVDD.n325 3.79678
R1039 AVDD.n252 AVDD.n246 3.79678
R1040 AVDD.n205 AVDD.n199 3.79678
R1041 AVDD.n1863 AVDD.n1862 3.74038
R1042 AVDD.n270 AVDD.n269 3.74038
R1043 AVDD.n1893 AVDD.n1887 3.73034
R1044 AVDD.n1844 AVDD.n1820 3.73034
R1045 AVDD.n338 AVDD.n314 3.73034
R1046 AVDD.n240 AVDD.n234 3.73034
R1047 AVDD.n1125 AVDD.t717 3.7109
R1048 AVDD.n1150 AVDD.n1149 3.68344
R1049 AVDD.n1214 AVDD.n1213 3.65594
R1050 AVDD.n2122 AVDD.n2121 3.65581
R1051 AVDD.n2125 AVDD.n2124 3.65581
R1052 AVDD.n2128 AVDD.n2127 3.65581
R1053 AVDD.n2131 AVDD.n2130 3.65581
R1054 AVDD.n57 AVDD.n56 3.65581
R1055 AVDD.n54 AVDD.n53 3.65581
R1056 AVDD.n51 AVDD.n50 3.65581
R1057 AVDD.n2063 AVDD.n2062 3.65581
R1058 AVDD.n2066 AVDD.n2065 3.65581
R1059 AVDD.n2069 AVDD.n2068 3.65581
R1060 AVDD.n2072 AVDD.n2071 3.65581
R1061 AVDD.n2060 AVDD.n2059 3.65581
R1062 AVDD.n2057 AVDD.n2056 3.65581
R1063 AVDD.n2054 AVDD.n2053 3.65581
R1064 AVDD.n1721 AVDD.n1720 3.65581
R1065 AVDD.n1718 AVDD.n1717 3.65581
R1066 AVDD.n1715 AVDD.n1714 3.65581
R1067 AVDD.n1712 AVDD.n1711 3.65581
R1068 AVDD.n84 AVDD.n83 3.65581
R1069 AVDD.n81 AVDD.n80 3.65581
R1070 AVDD.n78 AVDD.n77 3.65581
R1071 AVDD.n1674 AVDD.n1673 3.65581
R1072 AVDD.n1671 AVDD.n1670 3.65581
R1073 AVDD.n1668 AVDD.n1667 3.65581
R1074 AVDD.n1665 AVDD.n1664 3.65581
R1075 AVDD.n1661 AVDD.n1660 3.65581
R1076 AVDD.n1658 AVDD.n1657 3.65581
R1077 AVDD.n1655 AVDD.n1654 3.65581
R1078 AVDD.n1221 AVDD.n1220 3.6512
R1079 AVDD.n1208 AVDD.n1207 3.6512
R1080 AVDD.n1218 AVDD.n1217 3.6512
R1081 AVDD.n1211 AVDD.n1210 3.6512
R1082 AVDD.n2132 AVDD.n2131 3.64443
R1083 AVDD.n2073 AVDD.n2072 3.64443
R1084 AVDD.n1712 AVDD.n1709 3.64443
R1085 AVDD.n1665 AVDD.n1662 3.64443
R1086 AVDD.n969 AVDD.n968 3.6266
R1087 AVDD.n1014 AVDD.n1013 3.62041
R1088 AVDD.n1017 AVDD.n1016 3.62041
R1089 AVDD.n1021 AVDD.n1020 3.62041
R1090 AVDD.n1024 AVDD.n1023 3.62041
R1091 AVDD.n1027 AVDD.n1026 3.62041
R1092 AVDD.n728 AVDD.n727 3.61594
R1093 AVDD.n1968 AVDD.n1967 3.524
R1094 AVDD.n2089 AVDD.n2088 3.524
R1095 AVDD.n1991 AVDD.n1990 3.524
R1096 AVDD.n2027 AVDD.n2026 3.524
R1097 AVDD.n1553 AVDD.n1552 3.524
R1098 AVDD.n1683 AVDD.n1682 3.524
R1099 AVDD.n1600 AVDD.n1599 3.524
R1100 AVDD.n1633 AVDD.n1632 3.524
R1101 AVDD.n2077 AVDD.n2076 3.506
R1102 AVDD.n2015 AVDD.n2003 3.506
R1103 AVDD.n1689 AVDD.n1688 3.506
R1104 AVDD.n1639 AVDD.n1638 3.506
R1105 AVDD.n1727 AVDD.t138 3.20383
R1106 AVDD.n167 AVDD.t422 3.20383
R1107 AVDD.t384 AVDD.n168 3.20383
R1108 AVDD.n175 AVDD.t1076 3.20383
R1109 AVDD.t1108 AVDD.n176 3.20383
R1110 AVDD.t934 AVDD.n157 3.20383
R1111 AVDD.n2138 AVDD.t1208 3.20383
R1112 AVDD.n1740 AVDD.t1064 3.20383
R1113 AVDD.t1136 AVDD.n1741 3.20383
R1114 AVDD.n1748 AVDD.t418 3.20383
R1115 AVDD.t287 AVDD.n1749 3.20383
R1116 AVDD.t1168 AVDD.n1730 3.20383
R1117 AVDD.t104 AVDD.n1314 3.20383
R1118 AVDD.n1315 AVDD.t104 3.20383
R1119 AVDD.n1316 AVDD.t665 3.20383
R1120 AVDD.n1325 AVDD.t904 3.20383
R1121 AVDD.t527 AVDD.n1326 3.20383
R1122 AVDD.n1333 AVDD.t501 3.20383
R1123 AVDD.n1334 AVDD.t90 3.20383
R1124 AVDD.n1343 AVDD.t1098 3.20383
R1125 AVDD.t9 AVDD.n1344 3.20383
R1126 AVDD.n1345 AVDD.t9 3.20383
R1127 AVDD.t938 AVDD.n1350 3.20383
R1128 AVDD.n1351 AVDD.t938 3.20383
R1129 AVDD.n1352 AVDD.t1158 3.20383
R1130 AVDD.n1361 AVDD.t426 3.20383
R1131 AVDD.t1016 AVDD.n1362 3.20383
R1132 AVDD.n1369 AVDD.t6 3.20383
R1133 AVDD.n1370 AVDD.t594 3.20383
R1134 AVDD.n1379 AVDD.t1210 3.20383
R1135 AVDD.n1314 AVDD.t116 3.20383
R1136 AVDD.n1315 AVDD.t116 3.20383
R1137 AVDD.n1316 AVDD.t673 3.20383
R1138 AVDD.n1325 AVDD.t910 3.20383
R1139 AVDD.n1326 AVDD.t533 3.20383
R1140 AVDD.n1333 AVDD.t509 3.20383
R1141 AVDD.n1334 AVDD.t102 3.20383
R1142 AVDD.n1343 AVDD.t1104 3.20383
R1143 AVDD.n1344 AVDD.t25 3.20383
R1144 AVDD.n1345 AVDD.t25 3.20383
R1145 AVDD.n1350 AVDD.t942 3.20383
R1146 AVDD.n1351 AVDD.t942 3.20383
R1147 AVDD.n1352 AVDD.t1166 3.20383
R1148 AVDD.n1361 AVDD.t430 3.20383
R1149 AVDD.n1362 AVDD.t1020 3.20383
R1150 AVDD.n1369 AVDD.t11 3.20383
R1151 AVDD.n1370 AVDD.t600 3.20383
R1152 AVDD.n1379 AVDD.t1216 3.20383
R1153 AVDD.n1290 AVDD.t1246 3.20383
R1154 AVDD.t1246 AVDD.n1289 3.20383
R1155 AVDD.n1288 AVDD.t715 3.20383
R1156 AVDD.n1278 AVDD.t900 3.20383
R1157 AVDD.n1277 AVDD.t620 3.20383
R1158 AVDD.t239 AVDD.n1270 3.20383
R1159 AVDD.n1269 AVDD.t489 3.20383
R1160 AVDD.t206 AVDD.n32 3.20383
R1161 AVDD.n1949 AVDD.t819 3.20383
R1162 AVDD.n1940 AVDD.t996 3.20383
R1163 AVDD.n1939 AVDD.t732 3.20383
R1164 AVDD.t343 AVDD.n1932 3.20383
R1165 AVDD.n1931 AVDD.t586 3.20383
R1166 AVDD.t311 AVDD.n42 3.20383
R1167 AVDD.n2164 AVDD.t1112 3.20383
R1168 AVDD.n2173 AVDD.t988 3.20383
R1169 AVDD.t1024 AVDD.n2174 3.20383
R1170 AVDD.n1388 AVDD.t331 3.20383
R1171 AVDD.n1389 AVDD.t153 3.20383
R1172 AVDD.n1398 AVDD.t1056 3.20383
R1173 AVDD.n2164 AVDD.t466 3.20383
R1174 AVDD.n2173 AVDD.t341 3.20383
R1175 AVDD.n2174 AVDD.t376 3.20383
R1176 AVDD.n1388 AVDD.t964 3.20383
R1177 AVDD.n1389 AVDD.t813 3.20383
R1178 AVDD.n1398 AVDD.t412 3.20383
R1179 AVDD.n553 AVDD.t736 3.20383
R1180 AVDD.n543 AVDD.t699 3.20383
R1181 AVDD.n542 AVDD.t970 3.20383
R1182 AVDD.t382 AVDD.n535 3.20383
R1183 AVDD.n534 AVDD.t348 3.20383
R1184 AVDD.n524 AVDD.t1200 3.20383
R1185 AVDD.n523 AVDD.t150 3.20383
R1186 AVDD.t150 AVDD.n522 3.20383
R1187 AVDD.n553 AVDD.t1140 3.20383
R1188 AVDD.t1078 AVDD.n543 3.20383
R1189 AVDD.n542 AVDD.t60 3.20383
R1190 AVDD.n535 AVDD.t804 3.20383
R1191 AVDD.n534 AVDD.t758 3.20383
R1192 AVDD.t333 AVDD.n524 3.20383
R1193 AVDD.n523 AVDD.t570 3.20383
R1194 AVDD.n522 AVDD.t570 3.20383
R1195 AVDD.t558 AVDD.n12 3.20383
R1196 AVDD.n471 AVDD.t839 3.20383
R1197 AVDD.t796 AVDD.n472 3.20383
R1198 AVDD.n479 AVDD.t201 3.20383
R1199 AVDD.n480 AVDD.t227 3.20383
R1200 AVDD.n489 AVDD.t1280 3.20383
R1201 AVDD.t950 AVDD.n12 3.20383
R1202 AVDD.n471 AVDD.t1218 3.20383
R1203 AVDD.n472 AVDD.t1176 3.20383
R1204 AVDD.n479 AVDD.t612 3.20383
R1205 AVDD.n480 AVDD.t630 3.20383
R1206 AVDD.n489 AVDD.t434 3.20383
R1207 AVDD.n1465 AVDD.t454 3.20383
R1208 AVDD.n1474 AVDD.t762 3.20383
R1209 AVDD.t156 AVDD.n1475 3.20383
R1210 AVDD.t1146 AVDD.n665 3.20383
R1211 AVDD.n662 AVDD.t462 3.20383
R1212 AVDD.n652 AVDD.t244 3.20383
R1213 AVDD.n651 AVDD.t968 3.20383
R1214 AVDD.t968 AVDD.n650 3.20383
R1215 AVDD.n648 AVDD.t408 3.20383
R1216 AVDD.t408 AVDD.n647 3.20383
R1217 AVDD.n646 AVDD.t1148 3.20383
R1218 AVDD.n636 AVDD.t460 3.20383
R1219 AVDD.n635 AVDD.t859 3.20383
R1220 AVDD.t531 AVDD.n628 3.20383
R1221 AVDD.n627 AVDD.t1224 3.20383
R1222 AVDD.n617 AVDD.t821 3.20383
R1223 AVDD.n616 AVDD.t592 3.20383
R1224 AVDD.t592 AVDD.n615 3.20383
R1225 AVDD.n1465 AVDD.t464 3.20383
R1226 AVDD.n1474 AVDD.t770 3.20383
R1227 AVDD.n1475 AVDD.t160 3.20383
R1228 AVDD.n665 AVDD.t1152 3.20383
R1229 AVDD.n662 AVDD.t474 3.20383
R1230 AVDD.t250 AVDD.n652 3.20383
R1231 AVDD.n651 AVDD.t976 3.20383
R1232 AVDD.n650 AVDD.t976 3.20383
R1233 AVDD.n648 AVDD.t410 3.20383
R1234 AVDD.n647 AVDD.t410 3.20383
R1235 AVDD.n646 AVDD.t1156 3.20383
R1236 AVDD.t468 AVDD.n636 3.20383
R1237 AVDD.n635 AVDD.t861 3.20383
R1238 AVDD.n628 AVDD.t539 3.20383
R1239 AVDD.n627 AVDD.t1230 3.20383
R1240 AVDD.t829 AVDD.n617 3.20383
R1241 AVDD.n616 AVDD.t598 3.20383
R1242 AVDD.n615 AVDD.t598 3.20383
R1243 AVDD.n570 AVDD.t275 3.20383
R1244 AVDD.n579 AVDD.t218 3.20383
R1245 AVDD.t491 AVDD.n580 3.20383
R1246 AVDD.n587 AVDD.t1190 3.20383
R1247 AVDD.n588 AVDD.t1160 3.20383
R1248 AVDD.n597 AVDD.t750 3.20383
R1249 AVDD.t51 AVDD.n15 3.20383
R1250 AVDD.n430 AVDD.t360 3.20383
R1251 AVDD.t317 AVDD.n431 3.20383
R1252 AVDD.n438 AVDD.t1012 3.20383
R1253 AVDD.n439 AVDD.t1028 3.20383
R1254 AVDD.n448 AVDD.t873 3.20383
R1255 AVDD.n1506 AVDD.t242 3.20383
R1256 AVDD.n1515 AVDD.t193 3.20383
R1257 AVDD.t456 AVDD.n1516 3.20383
R1258 AVDD.n383 AVDD.t1172 3.20383
R1259 AVDD.n384 AVDD.t1128 3.20383
R1260 AVDD.n393 AVDD.t728 3.20383
R1261 AVDD.n394 AVDD.t952 3.20383
R1262 AVDD.t952 AVDD.n374 3.20383
R1263 AVDD.n1506 AVDD.t886 3.20383
R1264 AVDD.n1515 AVDD.t847 3.20383
R1265 AVDD.n1516 AVDD.t1092 3.20383
R1266 AVDD.n383 AVDD.t525 3.20383
R1267 AVDD.n384 AVDD.t483 3.20383
R1268 AVDD.n393 AVDD.t45 3.20383
R1269 AVDD.n394 AVDD.t309 3.20383
R1270 AVDD.t309 AVDD.n374 3.20383
R1271 AVDD.n1538 AVDD.t345 3.20383
R1272 AVDD.n1529 AVDD.t307 3.20383
R1273 AVDD.n1528 AVDD.t576 3.20383
R1274 AVDD.n351 AVDD.t1254 3.20383
R1275 AVDD.n352 AVDD.t1214 3.20383
R1276 AVDD.n361 AVDD.t827 3.20383
R1277 AVDD.n1438 AVDD.t23 3.20383
R1278 AVDD.n1428 AVDD.t339 3.20383
R1279 AVDD.n1427 AVDD.t299 3.20383
R1280 AVDD.t994 AVDD.n1420 3.20383
R1281 AVDD.n1419 AVDD.t1010 3.20383
R1282 AVDD.t845 AVDD.n109 3.20383
R1283 AVDD.n1438 AVDD.t693 3.20383
R1284 AVDD.t974 AVDD.n1428 3.20383
R1285 AVDD.n1427 AVDD.t928 3.20383
R1286 AVDD.n1420 AVDD.t352 3.20383
R1287 AVDD.n1419 AVDD.t369 3.20383
R1288 AVDD.t178 AVDD.n109 3.20383
R1289 AVDD.n768 AVDD.t922 3.20383
R1290 AVDD.n765 AVDD.t641 3.20383
R1291 AVDD.t273 AVDD.n761 3.20383
R1292 AVDD.n757 AVDD.t511 3.20383
R1293 AVDD.t229 AVDD.n939 3.20383
R1294 AVDD.n935 AVDD.t1250 3.20383
R1295 AVDD.t1250 AVDD.n934 3.20383
R1296 AVDD.n928 AVDD.t77 3.20383
R1297 AVDD.t77 AVDD.n927 3.20383
R1298 AVDD.n924 AVDD.t1154 3.20383
R1299 AVDD.t655 AVDD.n713 3.20383
R1300 AVDD.n714 AVDD.t655 3.20383
R1301 AVDD.t1204 AVDD.n770 3.20383
R1302 AVDD.n781 AVDD.t1252 3.20383
R1303 AVDD.n945 AVDD.t1044 3.20383
R1304 AVDD.t28 AVDD.n942 3.20383
R1305 AVDD.n938 AVDD.t687 3.20383
R1306 AVDD.n925 AVDD.t476 3.20383
R1307 AVDD.t616 AVDD.n906 3.20383
R1308 AVDD.n916 AVDD.t616 3.20383
R1309 AVDD.n1233 AVDD.t740 3.20383
R1310 AVDD.t1006 AVDD.n912 3.20383
R1311 AVDD.n911 AVDD.t1042 3.20383
R1312 AVDD.n2185 AVDD.t356 3.20383
R1313 AVDD.n2186 AVDD.t183 3.20383
R1314 AVDD.n2195 AVDD.t1074 3.20383
R1315 AVDD.n879 AVDD.t336 3.20383
R1316 AVDD.n869 AVDD.t196 3.20383
R1317 AVDD.n868 AVDD.t253 3.20383
R1318 AVDD.t835 AVDD.n861 3.20383
R1319 AVDD.n860 AVDD.t663 3.20383
R1320 AVDD.t295 AVDD.n13 3.20383
R1321 AVDD.n879 AVDD.t746 3.20383
R1322 AVDD.t602 AVDD.n869 3.20383
R1323 AVDD.n868 AVDD.t647 3.20383
R1324 AVDD.n861 AVDD.t1212 3.20383
R1325 AVDD.n860 AVDD.t1054 3.20383
R1326 AVDD.t683 AVDD.n13 3.20383
R1327 AVDD.t478 AVDD.n809 3.20383
R1328 AVDD.n810 AVDD.t478 3.20383
R1329 AVDD.n811 AVDD.t1198 3.20383
R1330 AVDD.n820 AVDD.t93 3.20383
R1331 AVDD.t1102 AVDD.n821 3.20383
R1332 AVDD.n828 AVDD.t734 3.20383
R1333 AVDD.n829 AVDD.t986 3.20383
R1334 AVDD.n838 AVDD.t709 3.20383
R1335 AVDD.n809 AVDD.t896 3.20383
R1336 AVDD.n810 AVDD.t896 3.20383
R1337 AVDD.n811 AVDD.t326 3.20383
R1338 AVDD.n820 AVDD.t507 3.20383
R1339 AVDD.n821 AVDD.t234 3.20383
R1340 AVDD.n828 AVDD.t1138 3.20383
R1341 AVDD.n829 AVDD.t83 3.20383
R1342 AVDD.n838 AVDD.t1088 3.20383
R1343 AVDD.n1095 AVDD.t811 3.20383
R1344 AVDD.n1086 AVDD.t876 3.20383
R1345 AVDD.n1085 AVDD.t639 3.20383
R1346 AVDD.t926 AVDD.n1078 3.20383
R1347 AVDD.n1077 AVDD.t283 3.20383
R1348 AVDD.n1068 AVDD.t40 3.20383
R1349 AVDD.n1290 AVDD.t622 3.20383
R1350 AVDD.n1289 AVDD.t622 3.20383
R1351 AVDD.n1288 AVDD.t34 3.20383
R1352 AVDD.t258 AVDD.n1278 3.20383
R1353 AVDD.n1277 AVDD.t1240 3.20383
R1354 AVDD.n1270 AVDD.t884 3.20383
R1355 AVDD.n1269 AVDD.t1114 3.20383
R1356 AVDD.t851 AVDD.n32 3.20383
R1357 AVDD.n1921 AVDD.n1920 3.00663
R1358 AVDD.n1853 AVDD.n1852 3.00663
R1359 AVDD.n341 AVDD.n154 3.00663
R1360 AVDD.n263 AVDD.n262 3.00663
R1361 AVDD.n1868 AVDD.n1865 2.7866
R1362 AVDD.n1873 AVDD.n1870 2.7866
R1363 AVDD.n1879 AVDD.n1876 2.7866
R1364 AVDD.n1885 AVDD.n1882 2.7866
R1365 AVDD.n1892 AVDD.n1889 2.7866
R1366 AVDD.n1898 AVDD.n1895 2.7866
R1367 AVDD.n1904 AVDD.n1901 2.7866
R1368 AVDD.n1910 AVDD.n1907 2.7866
R1369 AVDD.n1825 AVDD.n1822 2.7866
R1370 AVDD.n1830 AVDD.n1827 2.7866
R1371 AVDD.n1836 AVDD.n1833 2.7866
R1372 AVDD.n1842 AVDD.n1839 2.7866
R1373 AVDD.n1819 AVDD.n1816 2.7866
R1374 AVDD.n1813 AVDD.n1810 2.7866
R1375 AVDD.n1807 AVDD.n1804 2.7866
R1376 AVDD.n1801 AVDD.n1798 2.7866
R1377 AVDD.n319 AVDD.n316 2.7866
R1378 AVDD.n324 AVDD.n321 2.7866
R1379 AVDD.n330 AVDD.n327 2.7866
R1380 AVDD.n336 AVDD.n333 2.7866
R1381 AVDD.n313 AVDD.n310 2.7866
R1382 AVDD.n307 AVDD.n304 2.7866
R1383 AVDD.n301 AVDD.n298 2.7866
R1384 AVDD.n295 AVDD.n292 2.7866
R1385 AVDD.n193 AVDD.n190 2.7866
R1386 AVDD.n198 AVDD.n195 2.7866
R1387 AVDD.n204 AVDD.n201 2.7866
R1388 AVDD.n210 AVDD.n207 2.7866
R1389 AVDD.n239 AVDD.n236 2.7866
R1390 AVDD.n245 AVDD.n242 2.7866
R1391 AVDD.n251 AVDD.n248 2.7866
R1392 AVDD.n257 AVDD.n254 2.7866
R1393 AVDD.n2108 AVDD.n2106 2.73714
R1394 AVDD.n2010 AVDD.n2008 2.73714
R1395 AVDD.n1697 AVDD.n1695 2.73714
R1396 AVDD.n1588 AVDD.n1586 2.73714
R1397 AVDD.n1874 AVDD.n1868 2.73672
R1398 AVDD.n1831 AVDD.n1825 2.73672
R1399 AVDD.n325 AVDD.n319 2.73672
R1400 AVDD.n199 AVDD.n193 2.73672
R1401 AVDD.n1028 AVDD.n1027 2.60496
R1402 AVDD.n1208 AVDD.n1205 2.60386
R1403 AVDD.n1061 AVDD.n1060 2.6005
R1404 AVDD.n1064 AVDD.n1063 2.6005
R1405 AVDD.n1038 AVDD.n1037 2.6005
R1406 AVDD.n1035 AVDD.n1034 2.6005
R1407 AVDD.n1014 AVDD.n1011 2.59852
R1408 AVDD.n1222 AVDD.n1221 2.59742
R1409 AVDD.n2046 AVDD.n2043 2.59712
R1410 AVDD.n2008 AVDD.n2005 2.59712
R1411 AVDD.n2114 AVDD.n2111 2.59712
R1412 AVDD.n2106 AVDD.n2103 2.59712
R1413 AVDD.n1646 AVDD.n1643 2.59712
R1414 AVDD.n1586 AVDD.n1583 2.59712
R1415 AVDD.n1704 AVDD.n1701 2.59712
R1416 AVDD.n1695 AVDD.n1692 2.59712
R1417 AVDD.n1042 AVDD.t1276 2.5255
R1418 AVDD.n1044 AVDD.t920 2.5255
R1419 AVDD.n1047 AVDD.t543 2.5255
R1420 AVDD.n1047 AVDD.t888 2.5255
R1421 AVDD.n1051 AVDD.t808 2.5255
R1422 AVDD.n1051 AVDD.t1132 2.5255
R1423 AVDD.n1054 AVDD.t436 2.5255
R1424 AVDD.n1054 AVDD.t798 2.5255
R1425 AVDD.n1056 AVDD.t3 2.5255
R1426 AVDD.n1056 AVDD.t374 2.5255
R1427 AVDD.n1031 AVDD.t14 2.5255
R1428 AVDD.n1005 AVDD.t932 2.5255
R1429 AVDD.n1000 AVDD.t898 2.5255
R1430 AVDD.n1119 AVDD.t1150 2.5255
R1431 AVDD.n989 AVDD.t806 2.5255
R1432 AVDD.n1066 AVDD.t388 2.5255
R1433 AVDD.n1200 AVDD.n1199 2.46986
R1434 AVDD.n1132 AVDD.n1131 2.46873
R1435 AVDD.n1117 AVDD.n1116 2.46873
R1436 AVDD.n1099 AVDD.n1098 2.46198
R1437 AVDD.n1178 AVDD.n1177 2.46198
R1438 AVDD.n1182 AVDD.n1181 2.46086
R1439 AVDD.n2109 AVDD.n2108 2.46014
R1440 AVDD.n2048 AVDD.n2010 2.46014
R1441 AVDD.n1706 AVDD.n1697 2.46014
R1442 AVDD.n1641 AVDD.n1588 2.46014
R1443 AVDD.n1034 AVDD.t395 2.4505
R1444 AVDD.n1034 AVDD.t329 2.4505
R1445 AVDD.t1184 AVDD.n1038 2.4505
R1446 AVDD.n1038 AVDD.t395 2.4505
R1447 AVDD.n1064 AVDD.t742 2.4505
R1448 AVDD.t667 AVDD.n1064 2.4505
R1449 AVDD.n1060 AVDD.t265 2.4505
R1450 AVDD.n1060 AVDD.t742 2.4505
R1451 AVDD.n2046 AVDD.n2045 2.39107
R1452 AVDD.n2008 AVDD.n2007 2.39107
R1453 AVDD.n2114 AVDD.n2113 2.39107
R1454 AVDD.n2106 AVDD.n2105 2.39107
R1455 AVDD.n1646 AVDD.n1645 2.39107
R1456 AVDD.n1586 AVDD.n1585 2.39107
R1457 AVDD.n1704 AVDD.n1703 2.39107
R1458 AVDD.n1695 AVDD.n1694 2.39107
R1459 AVDD.n1789 AVDD.n1788 2.37568
R1460 AVDD.n1765 AVDD.n1764 2.37568
R1461 AVDD.n221 AVDD.n220 2.37568
R1462 AVDD.n278 AVDD.n277 2.37568
R1463 AVDD.n1176 AVDD.n1175 2.37449
R1464 AVDD.n1168 AVDD.n1167 2.37449
R1465 AVDD.n1160 AVDD.n1159 2.37449
R1466 AVDD.n1146 AVDD.n1145 2.37449
R1467 AVDD.n1138 AVDD.n1137 2.37449
R1468 AVDD.n2134 AVDD.n43 2.30165
R1469 AVDD.n1951 AVDD.n1950 2.30165
R1470 AVDD.n1723 AVDD.n70 2.30165
R1471 AVDD.n1540 AVDD.n1539 2.30165
R1472 AVDD.n1856 AVDD.n1773 2.24038
R1473 AVDD.n1782 AVDD.n1781 2.24038
R1474 AVDD.n289 AVDD.n288 2.24038
R1475 AVDD.n232 AVDD.n231 2.24038
R1476 AVDD.n1173 AVDD.n1172 2.21344
R1477 AVDD.n1165 AVDD.n1164 2.21344
R1478 AVDD.n1157 AVDD.n1156 2.21344
R1479 AVDD.n1143 AVDD.n1142 2.21344
R1480 AVDD.n1135 AVDD.n1134 2.21344
R1481 AVDD.n1868 AVDD.n1867 2.2016
R1482 AVDD.n1873 AVDD.n1872 2.2016
R1483 AVDD.n1879 AVDD.n1878 2.2016
R1484 AVDD.n1885 AVDD.n1884 2.2016
R1485 AVDD.n1892 AVDD.n1891 2.2016
R1486 AVDD.n1898 AVDD.n1897 2.2016
R1487 AVDD.n1904 AVDD.n1903 2.2016
R1488 AVDD.n1910 AVDD.n1909 2.2016
R1489 AVDD.n1825 AVDD.n1824 2.2016
R1490 AVDD.n1830 AVDD.n1829 2.2016
R1491 AVDD.n1836 AVDD.n1835 2.2016
R1492 AVDD.n1842 AVDD.n1841 2.2016
R1493 AVDD.n1819 AVDD.n1818 2.2016
R1494 AVDD.n1813 AVDD.n1812 2.2016
R1495 AVDD.n1807 AVDD.n1806 2.2016
R1496 AVDD.n1801 AVDD.n1800 2.2016
R1497 AVDD.n319 AVDD.n318 2.2016
R1498 AVDD.n324 AVDD.n323 2.2016
R1499 AVDD.n330 AVDD.n329 2.2016
R1500 AVDD.n336 AVDD.n335 2.2016
R1501 AVDD.n313 AVDD.n312 2.2016
R1502 AVDD.n307 AVDD.n306 2.2016
R1503 AVDD.n301 AVDD.n300 2.2016
R1504 AVDD.n295 AVDD.n294 2.2016
R1505 AVDD.n193 AVDD.n192 2.2016
R1506 AVDD.n198 AVDD.n197 2.2016
R1507 AVDD.n204 AVDD.n203 2.2016
R1508 AVDD.n210 AVDD.n209 2.2016
R1509 AVDD.n239 AVDD.n238 2.2016
R1510 AVDD.n245 AVDD.n244 2.2016
R1511 AVDD.n251 AVDD.n250 2.2016
R1512 AVDD.n257 AVDD.n256 2.2016
R1513 AVDD.n2039 AVDD.n2038 2.18645
R1514 AVDD.n1650 AVDD.n1581 2.18645
R1515 AVDD.n2098 AVDD.n2097 2.18502
R1516 AVDD.n2092 AVDD.n2091 2.18502
R1517 AVDD.n2086 AVDD.n2085 2.18502
R1518 AVDD.n2080 AVDD.n2079 2.18502
R1519 AVDD.n1977 AVDD.n1976 2.18502
R1520 AVDD.n1971 AVDD.n1970 2.18502
R1521 AVDD.n1965 AVDD.n1964 2.18502
R1522 AVDD.n2036 AVDD.n2035 2.18502
R1523 AVDD.n2030 AVDD.n2029 2.18502
R1524 AVDD.n2024 AVDD.n2023 2.18502
R1525 AVDD.n2018 AVDD.n2017 2.18502
R1526 AVDD.n2000 AVDD.n1999 2.18502
R1527 AVDD.n1994 AVDD.n1993 2.18502
R1528 AVDD.n1988 AVDD.n1987 2.18502
R1529 AVDD.n1580 AVDD.n1579 2.18502
R1530 AVDD.n1576 AVDD.n1575 2.18502
R1531 AVDD.n1572 AVDD.n1571 2.18502
R1532 AVDD.n1568 AVDD.n1567 2.18502
R1533 AVDD.n1562 AVDD.n1561 2.18502
R1534 AVDD.n1556 AVDD.n1555 2.18502
R1535 AVDD.n1550 AVDD.n1549 2.18502
R1536 AVDD.n1627 AVDD.n1626 2.18502
R1537 AVDD.n1623 AVDD.n1622 2.18502
R1538 AVDD.n1619 AVDD.n1618 2.18502
R1539 AVDD.n1615 AVDD.n1614 2.18502
R1540 AVDD.n1609 AVDD.n1608 2.18502
R1541 AVDD.n1603 AVDD.n1602 2.18502
R1542 AVDD.n1597 AVDD.n1596 2.18502
R1543 AVDD.n981 AVDD.n980 2.1566
R1544 AVDD.n977 AVDD.n976 2.1566
R1545 AVDD.n973 AVDD.n972 2.1566
R1546 AVDD.n966 AVDD.n965 2.1566
R1547 AVDD.n962 AVDD.n961 2.1566
R1548 AVDD.n740 AVDD.n739 2.14594
R1549 AVDD.n736 AVDD.n735 2.14594
R1550 AVDD.n732 AVDD.n731 2.14594
R1551 AVDD.n725 AVDD.n724 2.14594
R1552 AVDD.n721 AVDD.n720 2.14594
R1553 AVDD.n2049 AVDD.n2003 2.0852
R1554 AVDD.n1845 AVDD.n1782 2.0852
R1555 AVDD.n1640 AVDD.n1639 2.0852
R1556 AVDD.n233 AVDD.n232 2.0852
R1557 AVDD.n2122 AVDD.n2119 1.73609
R1558 AVDD.n2063 AVDD.n1952 1.73609
R1559 AVDD.n1722 AVDD.n1721 1.73609
R1560 AVDD.n1675 AVDD.n1674 1.73609
R1561 AVDD.n1925 AVDD.n1924 1.73383
R1562 AVDD.n1927 AVDD.n1926 1.73383
R1563 AVDD.n1930 AVDD.n1929 1.73383
R1564 AVDD.n1934 AVDD.n1933 1.73383
R1565 AVDD.n1938 AVDD.n1937 1.73383
R1566 AVDD.n1943 AVDD.n1942 1.73383
R1567 AVDD.n1945 AVDD.n1944 1.73383
R1568 AVDD.n1948 AVDD.n1947 1.73383
R1569 AVDD.n1396 AVDD.n1381 1.73383
R1570 AVDD.n1394 AVDD.n1382 1.73383
R1571 AVDD.n1391 AVDD.n1384 1.73383
R1572 AVDD.n1385 AVDD.n24 1.73383
R1573 AVDD.n2176 AVDD.n25 1.73383
R1574 AVDD.n2171 AVDD.n28 1.73383
R1575 AVDD.n2169 AVDD.n29 1.73383
R1576 AVDD.n2166 AVDD.n31 1.73383
R1577 AVDD.n1397 AVDD.n1396 1.73383
R1578 AVDD.n1394 AVDD.n1393 1.73383
R1579 AVDD.n1392 AVDD.n1391 1.73383
R1580 AVDD.n1387 AVDD.n24 1.73383
R1581 AVDD.n2176 AVDD.n2175 1.73383
R1582 AVDD.n2172 AVDD.n2171 1.73383
R1583 AVDD.n2169 AVDD.n2168 1.73383
R1584 AVDD.n2167 AVDD.n2166 1.73383
R1585 AVDD.n487 AVDD.n450 1.73383
R1586 AVDD.n485 AVDD.n451 1.73383
R1587 AVDD.n482 AVDD.n453 1.73383
R1588 AVDD.n477 AVDD.n455 1.73383
R1589 AVDD.n474 AVDD.n456 1.73383
R1590 AVDD.n469 AVDD.n459 1.73383
R1591 AVDD.n467 AVDD.n460 1.73383
R1592 AVDD.n464 AVDD.n462 1.73383
R1593 AVDD.n488 AVDD.n487 1.73383
R1594 AVDD.n485 AVDD.n484 1.73383
R1595 AVDD.n483 AVDD.n482 1.73383
R1596 AVDD.n478 AVDD.n477 1.73383
R1597 AVDD.n474 AVDD.n473 1.73383
R1598 AVDD.n470 AVDD.n469 1.73383
R1599 AVDD.n467 AVDD.n466 1.73383
R1600 AVDD.n465 AVDD.n464 1.73383
R1601 AVDD.n447 AVDD.n446 1.73383
R1602 AVDD.n444 AVDD.n443 1.73383
R1603 AVDD.n442 AVDD.n441 1.73383
R1604 AVDD.n437 AVDD.n436 1.73383
R1605 AVDD.n433 AVDD.n432 1.73383
R1606 AVDD.n429 AVDD.n428 1.73383
R1607 AVDD.n426 AVDD.n425 1.73383
R1608 AVDD.n424 AVDD.n423 1.73383
R1609 AVDD.n596 AVDD.n595 1.73383
R1610 AVDD.n593 AVDD.n592 1.73383
R1611 AVDD.n591 AVDD.n590 1.73383
R1612 AVDD.n586 AVDD.n585 1.73383
R1613 AVDD.n582 AVDD.n581 1.73383
R1614 AVDD.n578 AVDD.n577 1.73383
R1615 AVDD.n575 AVDD.n574 1.73383
R1616 AVDD.n573 AVDD.n572 1.73383
R1617 AVDD.n360 AVDD.n359 1.73383
R1618 AVDD.n357 AVDD.n356 1.73383
R1619 AVDD.n355 AVDD.n354 1.73383
R1620 AVDD.n350 AVDD.n90 1.73383
R1621 AVDD.n1527 AVDD.n1526 1.73383
R1622 AVDD.n1532 AVDD.n1531 1.73383
R1623 AVDD.n1534 AVDD.n1533 1.73383
R1624 AVDD.n1537 AVDD.n1536 1.73383
R1625 AVDD.n1411 AVDD.n1410 1.73383
R1626 AVDD.n1415 AVDD.n1414 1.73383
R1627 AVDD.n1417 AVDD.n1416 1.73383
R1628 AVDD.n1423 AVDD.n1422 1.73383
R1629 AVDD.n1425 AVDD.n1424 1.73383
R1630 AVDD.n1430 AVDD.n1429 1.73383
R1631 AVDD.n1434 AVDD.n1433 1.73383
R1632 AVDD.n1436 AVDD.n1435 1.73383
R1633 AVDD.n1412 AVDD.n1411 1.73383
R1634 AVDD.n1414 AVDD.n1413 1.73383
R1635 AVDD.n1418 AVDD.n1417 1.73383
R1636 AVDD.n1422 AVDD.n1421 1.73383
R1637 AVDD.n1426 AVDD.n1425 1.73383
R1638 AVDD.n1431 AVDD.n1430 1.73383
R1639 AVDD.n1433 AVDD.n1432 1.73383
R1640 AVDD.n1437 AVDD.n1436 1.73383
R1641 AVDD.n391 AVDD.n376 1.73383
R1642 AVDD.n389 AVDD.n377 1.73383
R1643 AVDD.n386 AVDD.n379 1.73383
R1644 AVDD.n380 AVDD.n101 1.73383
R1645 AVDD.n1518 AVDD.n102 1.73383
R1646 AVDD.n1513 AVDD.n105 1.73383
R1647 AVDD.n1511 AVDD.n106 1.73383
R1648 AVDD.n1508 AVDD.n108 1.73383
R1649 AVDD.n392 AVDD.n391 1.73383
R1650 AVDD.n389 AVDD.n388 1.73383
R1651 AVDD.n387 AVDD.n386 1.73383
R1652 AVDD.n382 AVDD.n101 1.73383
R1653 AVDD.n1518 AVDD.n1517 1.73383
R1654 AVDD.n1514 AVDD.n1513 1.73383
R1655 AVDD.n1511 AVDD.n1510 1.73383
R1656 AVDD.n1509 AVDD.n1508 1.73383
R1657 AVDD.n619 AVDD.n618 1.73383
R1658 AVDD.n623 AVDD.n622 1.73383
R1659 AVDD.n625 AVDD.n624 1.73383
R1660 AVDD.n631 AVDD.n630 1.73383
R1661 AVDD.n633 AVDD.n632 1.73383
R1662 AVDD.n638 AVDD.n637 1.73383
R1663 AVDD.n642 AVDD.n641 1.73383
R1664 AVDD.n644 AVDD.n643 1.73383
R1665 AVDD.n654 AVDD.n653 1.73383
R1666 AVDD.n658 AVDD.n657 1.73383
R1667 AVDD.n660 AVDD.n659 1.73383
R1668 AVDD.n663 AVDD.n122 1.73383
R1669 AVDD.n1477 AVDD.n123 1.73383
R1670 AVDD.n1472 AVDD.n668 1.73383
R1671 AVDD.n1470 AVDD.n669 1.73383
R1672 AVDD.n1467 AVDD.n671 1.73383
R1673 AVDD.n620 AVDD.n619 1.73383
R1674 AVDD.n622 AVDD.n621 1.73383
R1675 AVDD.n626 AVDD.n625 1.73383
R1676 AVDD.n630 AVDD.n629 1.73383
R1677 AVDD.n634 AVDD.n633 1.73383
R1678 AVDD.n639 AVDD.n638 1.73383
R1679 AVDD.n641 AVDD.n640 1.73383
R1680 AVDD.n645 AVDD.n644 1.73383
R1681 AVDD.n655 AVDD.n654 1.73383
R1682 AVDD.n657 AVDD.n656 1.73383
R1683 AVDD.n661 AVDD.n660 1.73383
R1684 AVDD.n666 AVDD.n122 1.73383
R1685 AVDD.n1477 AVDD.n1476 1.73383
R1686 AVDD.n1473 AVDD.n1472 1.73383
R1687 AVDD.n1470 AVDD.n1469 1.73383
R1688 AVDD.n1468 AVDD.n1467 1.73383
R1689 AVDD.n526 AVDD.n525 1.73383
R1690 AVDD.n530 AVDD.n529 1.73383
R1691 AVDD.n532 AVDD.n531 1.73383
R1692 AVDD.n538 AVDD.n537 1.73383
R1693 AVDD.n540 AVDD.n539 1.73383
R1694 AVDD.n545 AVDD.n544 1.73383
R1695 AVDD.n549 AVDD.n548 1.73383
R1696 AVDD.n551 AVDD.n550 1.73383
R1697 AVDD.n527 AVDD.n526 1.73383
R1698 AVDD.n529 AVDD.n528 1.73383
R1699 AVDD.n533 AVDD.n532 1.73383
R1700 AVDD.n537 AVDD.n536 1.73383
R1701 AVDD.n541 AVDD.n540 1.73383
R1702 AVDD.n546 AVDD.n545 1.73383
R1703 AVDD.n548 AVDD.n547 1.73383
R1704 AVDD.n552 AVDD.n551 1.73383
R1705 AVDD.n1232 AVDD.n1231 1.73383
R1706 AVDD.n2194 AVDD.n2193 1.73383
R1707 AVDD.n2191 AVDD.n2190 1.73383
R1708 AVDD.n2189 AVDD.n2188 1.73383
R1709 AVDD.n2184 AVDD.n2183 1.73383
R1710 AVDD.n910 AVDD.n909 1.73383
R1711 AVDD.n914 AVDD.n913 1.73383
R1712 AVDD.n919 AVDD.n918 1.73383
R1713 AVDD.n836 AVDD.n788 1.73383
R1714 AVDD.n834 AVDD.n789 1.73383
R1715 AVDD.n831 AVDD.n791 1.73383
R1716 AVDD.n826 AVDD.n793 1.73383
R1717 AVDD.n823 AVDD.n794 1.73383
R1718 AVDD.n818 AVDD.n797 1.73383
R1719 AVDD.n816 AVDD.n798 1.73383
R1720 AVDD.n813 AVDD.n800 1.73383
R1721 AVDD.n837 AVDD.n836 1.73383
R1722 AVDD.n834 AVDD.n833 1.73383
R1723 AVDD.n832 AVDD.n831 1.73383
R1724 AVDD.n827 AVDD.n826 1.73383
R1725 AVDD.n823 AVDD.n822 1.73383
R1726 AVDD.n819 AVDD.n818 1.73383
R1727 AVDD.n816 AVDD.n815 1.73383
R1728 AVDD.n814 AVDD.n813 1.73383
R1729 AVDD.n852 AVDD.n851 1.73383
R1730 AVDD.n856 AVDD.n855 1.73383
R1731 AVDD.n858 AVDD.n857 1.73383
R1732 AVDD.n864 AVDD.n863 1.73383
R1733 AVDD.n866 AVDD.n865 1.73383
R1734 AVDD.n871 AVDD.n870 1.73383
R1735 AVDD.n875 AVDD.n874 1.73383
R1736 AVDD.n877 AVDD.n876 1.73383
R1737 AVDD.n853 AVDD.n852 1.73383
R1738 AVDD.n855 AVDD.n854 1.73383
R1739 AVDD.n859 AVDD.n858 1.73383
R1740 AVDD.n863 AVDD.n862 1.73383
R1741 AVDD.n867 AVDD.n866 1.73383
R1742 AVDD.n872 AVDD.n871 1.73383
R1743 AVDD.n874 AVDD.n873 1.73383
R1744 AVDD.n878 AVDD.n877 1.73383
R1745 AVDD.n1071 AVDD.n1070 1.73383
R1746 AVDD.n1073 AVDD.n1072 1.73383
R1747 AVDD.n1076 AVDD.n1075 1.73383
R1748 AVDD.n1080 AVDD.n1079 1.73383
R1749 AVDD.n1084 AVDD.n1083 1.73383
R1750 AVDD.n1089 AVDD.n1088 1.73383
R1751 AVDD.n1091 AVDD.n1090 1.73383
R1752 AVDD.n1094 AVDD.n1093 1.73383
R1753 AVDD.n930 AVDD.n929 1.73383
R1754 AVDD.n932 AVDD.n931 1.73383
R1755 AVDD.n937 AVDD.n936 1.73383
R1756 AVDD.n943 AVDD.n753 1.73383
R1757 AVDD.n944 AVDD.n756 1.73383
R1758 AVDD.n780 AVDD.n779 1.73383
R1759 AVDD.n766 AVDD.n764 1.73383
R1760 AVDD.n772 AVDD.n771 1.73383
R1761 AVDD.n923 AVDD.n922 1.73383
R1762 AVDD.n941 AVDD.n940 1.73383
R1763 AVDD.n951 AVDD.n950 1.73383
R1764 AVDD.n949 AVDD.n948 1.73383
R1765 AVDD.n778 AVDD.n777 1.73383
R1766 AVDD.n776 AVDD.n775 1.73383
R1767 AVDD.n1227 AVDD.n1226 1.73383
R1768 AVDD.n1229 AVDD.n1228 1.73383
R1769 AVDD.n1261 AVDD.n1260 1.73383
R1770 AVDD.n1265 AVDD.n1264 1.73383
R1771 AVDD.n1267 AVDD.n1266 1.73383
R1772 AVDD.n1273 AVDD.n1272 1.73383
R1773 AVDD.n1275 AVDD.n1274 1.73383
R1774 AVDD.n1280 AVDD.n1279 1.73383
R1775 AVDD.n1284 AVDD.n1283 1.73383
R1776 AVDD.n1286 AVDD.n1285 1.73383
R1777 AVDD.n1262 AVDD.n1261 1.73383
R1778 AVDD.n1264 AVDD.n1263 1.73383
R1779 AVDD.n1268 AVDD.n1267 1.73383
R1780 AVDD.n1272 AVDD.n1271 1.73383
R1781 AVDD.n1276 AVDD.n1275 1.73383
R1782 AVDD.n1281 AVDD.n1280 1.73383
R1783 AVDD.n1283 AVDD.n1282 1.73383
R1784 AVDD.n1287 AVDD.n1286 1.73383
R1785 AVDD.n1377 AVDD.n673 1.73383
R1786 AVDD.n1375 AVDD.n674 1.73383
R1787 AVDD.n1372 AVDD.n676 1.73383
R1788 AVDD.n1367 AVDD.n678 1.73383
R1789 AVDD.n1364 AVDD.n679 1.73383
R1790 AVDD.n1359 AVDD.n682 1.73383
R1791 AVDD.n1357 AVDD.n683 1.73383
R1792 AVDD.n1354 AVDD.n685 1.73383
R1793 AVDD.n1341 AVDD.n690 1.73383
R1794 AVDD.n1339 AVDD.n691 1.73383
R1795 AVDD.n1336 AVDD.n693 1.73383
R1796 AVDD.n1331 AVDD.n695 1.73383
R1797 AVDD.n1328 AVDD.n697 1.73383
R1798 AVDD.n1323 AVDD.n700 1.73383
R1799 AVDD.n1321 AVDD.n701 1.73383
R1800 AVDD.n1318 AVDD.n703 1.73383
R1801 AVDD.n1378 AVDD.n1377 1.73383
R1802 AVDD.n1375 AVDD.n1374 1.73383
R1803 AVDD.n1373 AVDD.n1372 1.73383
R1804 AVDD.n1368 AVDD.n1367 1.73383
R1805 AVDD.n1364 AVDD.n1363 1.73383
R1806 AVDD.n1360 AVDD.n1359 1.73383
R1807 AVDD.n1357 AVDD.n1356 1.73383
R1808 AVDD.n1355 AVDD.n1354 1.73383
R1809 AVDD.n1342 AVDD.n1341 1.73383
R1810 AVDD.n1339 AVDD.n1338 1.73383
R1811 AVDD.n1337 AVDD.n1336 1.73383
R1812 AVDD.n1332 AVDD.n1331 1.73383
R1813 AVDD.n1328 AVDD.n1327 1.73383
R1814 AVDD.n1324 AVDD.n1323 1.73383
R1815 AVDD.n1321 AVDD.n1320 1.73383
R1816 AVDD.n1319 AVDD.n1318 1.73383
R1817 AVDD.n1756 AVDD.n1755 1.73383
R1818 AVDD.n1754 AVDD.n1753 1.73383
R1819 AVDD.n1751 AVDD.n1750 1.73383
R1820 AVDD.n1747 AVDD.n1746 1.73383
R1821 AVDD.n1743 AVDD.n1742 1.73383
R1822 AVDD.n1739 AVDD.n1738 1.73383
R1823 AVDD.n1736 AVDD.n1735 1.73383
R1824 AVDD.n2137 AVDD.n2136 1.73383
R1825 AVDD.n183 AVDD.n182 1.73383
R1826 AVDD.n181 AVDD.n180 1.73383
R1827 AVDD.n178 AVDD.n177 1.73383
R1828 AVDD.n174 AVDD.n173 1.73383
R1829 AVDD.n170 AVDD.n169 1.73383
R1830 AVDD.n166 AVDD.n165 1.73383
R1831 AVDD.n163 AVDD.n162 1.73383
R1832 AVDD.n1726 AVDD.n1725 1.73383
R1833 AVDD.n1913 AVDD.n1757 1.69136
R1834 AVDD.n1923 AVDD.n1922 1.69136
R1835 AVDD.n340 AVDD.n184 1.69136
R1836 AVDD.n347 AVDD.n346 1.69136
R1837 AVDD.n1912 AVDD.n1911 1.65018
R1838 AVDD.n1802 AVDD.n1796 1.65018
R1839 AVDD.n296 AVDD.n151 1.65018
R1840 AVDD.n259 AVDD.n258 1.65018
R1841 AVDD.n1728 AVDD.t432 1.60217
R1842 AVDD.n2225 AVDD.t954 1.60217
R1843 AVDD.n2222 AVDD.t855 1.60217
R1844 AVDD.n2 AVDD.t924 1.60217
R1845 AVDD.n1441 AVDD.t1106 1.60217
R1846 AVDD.n1443 AVDD.t350 1.60217
R1847 AVDD.n1728 AVDD.t1188 1.60217
R1848 AVDD.n2225 AVDD.t416 1.60217
R1849 AVDD.n2222 AVDD.t321 1.60217
R1850 AVDD.n2 AVDD.t392 1.60217
R1851 AVDD.n1441 AVDD.t588 1.60217
R1852 AVDD.n1443 AVDD.t1084 1.60217
R1853 AVDD.n1445 AVDD.t982 1.60217
R1854 AVDD.n1447 AVDD.t208 1.60217
R1855 AVDD.n1450 AVDD.t71 1.60217
R1856 AVDD.n1453 AVDD.t212 1.60217
R1857 AVDD.n1456 AVDD.t73 1.60217
R1858 AVDD.n1458 AVDD.t677 1.60217
R1859 AVDD.n1445 AVDD.t442 1.60217
R1860 AVDD.n1447 AVDD.t960 1.60217
R1861 AVDD.n1450 AVDD.t867 1.60217
R1862 AVDD.n1453 AVDD.t222 1.60217
R1863 AVDD.n1456 AVDD.t114 1.60217
R1864 AVDD.n1458 AVDD.t695 1.60217
R1865 AVDD.n1463 AVDD.t681 1.60217
R1866 AVDD.n1461 AVDD.t1178 1.60217
R1867 AVDD.n10 AVDD.t1060 1.60217
R1868 AVDD.n2216 AVDD.t1066 1.60217
R1869 AVDD.n2213 AVDD.t760 1.60217
R1870 AVDD.n2211 AVDD.t849 1.60217
R1871 AVDD.n1463 AVDD.t703 1.60217
R1872 AVDD.n1461 AVDD.t1192 1.60217
R1873 AVDD.n10 AVDD.t1070 1.60217
R1874 AVDD.n2216 AVDD.t1090 1.60217
R1875 AVDD.n2213 AVDD.t262 1.60217
R1876 AVDD.n2211 AVDD.t315 1.60217
R1877 AVDD.n2209 AVDD.t1226 1.60217
R1878 AVDD.n2207 AVDD.t669 1.60217
R1879 AVDD.n2204 AVDD.t794 1.60217
R1880 AVDD.n2202 AVDD.t782 1.60217
R1881 AVDD.n2199 AVDD.t890 1.60217
R1882 AVDD.n2197 AVDD.t371 1.60217
R1883 AVDD.n2209 AVDD.t726 1.60217
R1884 AVDD.n2207 AVDD.t128 1.60217
R1885 AVDD.n2204 AVDD.t267 1.60217
R1886 AVDD.n2202 AVDD.t248 1.60217
R1887 AVDD.n2199 AVDD.t354 1.60217
R1888 AVDD.n2197 AVDD.t1120 1.60217
R1889 AVDD.n2140 AVDD.t47 1.60217
R1890 AVDD.n2142 AVDD.t584 1.60217
R1891 AVDD.n2145 AVDD.t452 1.60217
R1892 AVDD.n2151 AVDD.t551 1.60217
R1893 AVDD.n2148 AVDD.t752 1.60217
R1894 AVDD.n33 AVDD.t1236 1.60217
R1895 AVDD.n2140 AVDD.t168 1.60217
R1896 AVDD.n2142 AVDD.t691 1.60217
R1897 AVDD.n2145 AVDD.t578 1.60217
R1898 AVDD.n2151 AVDD.t651 1.60217
R1899 AVDD.n2148 AVDD.t863 1.60217
R1900 AVDD.n33 AVDD.t49 1.60217
R1901 AVDD.n2162 AVDD.t606 1.60217
R1902 AVDD.n2160 AVDD.t1100 1.60217
R1903 AVDD.n2157 AVDD.t1000 1.60217
R1904 AVDD.n34 AVDD.t882 1.60217
R1905 AVDD.n1348 AVDD.t774 1.60217
R1906 AVDD.n2162 AVDD.t720 1.60217
R1907 AVDD.n2160 AVDD.t1206 1.60217
R1908 AVDD.n2157 AVDD.t1096 1.60217
R1909 AVDD.n34 AVDD.t458 1.60217
R1910 AVDD.n1348 AVDD.t358 1.60217
R1911 AVDD.n1312 AVDD.t626 1.60217
R1912 AVDD.n1309 AVDD.t515 1.60217
R1913 AVDD.n706 AVDD.t521 1.60217
R1914 AVDD.n807 AVDD.t1196 1.60217
R1915 AVDD.n1298 AVDD.t1130 1.60217
R1916 AVDD.n1295 AVDD.t1014 1.60217
R1917 AVDD.n1293 AVDD.t936 1.60217
R1918 AVDD.n705 AVDD.t833 1.60217
R1919 AVDD.n60 AVDD.t63 1.60217
R1920 AVDD.n1243 AVDD.t596 1.60217
R1921 AVDD.n1246 AVDD.t487 1.60217
R1922 AVDD.n1303 AVDD.t564 1.60217
R1923 AVDD.n1300 AVDD.t776 1.60217
R1924 AVDD.n520 AVDD.t1256 1.60217
R1925 AVDD.n408 AVDD.t100 1.60217
R1926 AVDD.n603 AVDD.t68 1.60217
R1927 AVDD.n600 AVDD.t203 1.60217
R1928 AVDD.n598 AVDD.t980 1.60217
R1929 AVDD.n613 AVDD.t1094 1.60217
R1930 AVDD.n610 AVDD.t998 1.60217
R1931 AVDD.n514 AVDD.t1004 1.60217
R1932 AVDD.n517 AVDD.t636 1.60217
R1933 AVDD.n133 AVDD.t198 1.60217
R1934 AVDD.n492 AVDD.t57 1.60217
R1935 AVDD.n495 AVDD.t75 1.60217
R1936 AVDD.n498 AVDD.t547 1.60217
R1937 AVDD.n500 AVDD.t604 1.60217
R1938 AVDD.n133 AVDD.t930 1.60217
R1939 AVDD.n492 AVDD.t825 1.60217
R1940 AVDD.n495 AVDD.t843 1.60217
R1941 AVDD.n498 AVDD.t831 1.60217
R1942 AVDD.n500 AVDD.t162 1.60217
R1943 AVDD.n555 AVDD.t1002 1.60217
R1944 AVDD.n557 AVDD.t420 1.60217
R1945 AVDD.n560 AVDD.t545 1.60217
R1946 AVDD.n563 AVDD.t529 1.60217
R1947 AVDD.n566 AVDD.t634 1.60217
R1948 AVDD.n568 AVDD.t126 1.60217
R1949 AVDD.n555 AVDD.t582 1.60217
R1950 AVDD.n557 AVDD.t1258 1.60217
R1951 AVDD.n560 AVDD.t108 1.60217
R1952 AVDD.n563 AVDD.t80 1.60217
R1953 AVDD.n566 AVDD.t214 1.60217
R1954 AVDD.n568 AVDD.t990 1.60217
R1955 AVDD.n1483 AVDD.t210 1.60217
R1956 AVDD.n1485 AVDD.t730 1.60217
R1957 AVDD.n1488 AVDD.t608 1.60217
R1958 AVDD.n1493 AVDD.t685 1.60217
R1959 AVDD.n1490 AVDD.t894 1.60217
R1960 AVDD.n110 AVDD.t95 1.60217
R1961 AVDD.n1483 AVDD.t1050 1.60217
R1962 AVDD.n1485 AVDD.t301 1.60217
R1963 AVDD.n1488 AVDD.t166 1.60217
R1964 AVDD.n1493 AVDD.t271 1.60217
R1965 AVDD.n1490 AVDD.t440 1.60217
R1966 AVDD.n110 AVDD.t958 1.60217
R1967 AVDD.n1504 AVDD.t754 1.60217
R1968 AVDD.n1502 AVDD.t1238 1.60217
R1969 AVDD.n1499 AVDD.t1144 1.60217
R1970 AVDD.n111 AVDD.t499 1.60217
R1971 AVDD.n132 AVDD.t390 1.60217
R1972 AVDD.n1504 AVDD.t319 1.60217
R1973 AVDD.n1502 AVDD.t837 1.60217
R1974 AVDD.n1499 AVDD.t722 1.60217
R1975 AVDD.n111 AVDD.t1220 1.60217
R1976 AVDD.n132 AVDD.t1116 1.60217
R1977 AVDD.n397 AVDD.t823 1.60217
R1978 AVDD.n400 AVDD.t711 1.60217
R1979 AVDD.n403 AVDD.t124 1.60217
R1980 AVDD.n406 AVDD.t1272 1.60217
R1981 AVDD.n362 AVDD.t1038 1.60217
R1982 AVDD.n364 AVDD.t297 1.60217
R1983 AVDD.n367 AVDD.t158 1.60217
R1984 AVDD.n370 AVDD.t260 1.60217
R1985 AVDD.n373 AVDD.t428 1.60217
R1986 AVDD.n752 AVDD.t1080 1.60217
R1987 AVDD.n1003 AVDD.t659 1.60217
R1988 AVDD.n1120 AVDD.t784 1.60217
R1989 AVDD.n992 AVDD.t190 1.60217
R1990 AVDD.n1204 AVDD.t946 1.60217
R1991 AVDD.n1201 AVDD.t131 1.60217
R1992 AVDD.n751 AVDD.t679 1.60217
R1993 AVDD.n804 AVDD.t313 1.60217
R1994 AVDD.n711 AVDD.t414 1.60217
R1995 AVDD.n1239 AVDD.t406 1.60217
R1996 AVDD.n1236 AVDD.t517 1.60217
R1997 AVDD.n1234 AVDD.t1262 1.60217
R1998 AVDD.n687 AVDD.t566 1.60217
R1999 AVDD.n882 AVDD.t438 1.60217
R2000 AVDD.n885 AVDD.t450 1.60217
R2001 AVDD.n888 AVDD.t1018 1.60217
R2002 AVDD.n890 AVDD.t448 1.60217
R2003 AVDD.n687 AVDD.t143 1.60217
R2004 AVDD.n882 AVDD.t17 1.60217
R2005 AVDD.n885 AVDD.t42 1.60217
R2006 AVDD.n888 AVDD.t701 1.60217
R2007 AVDD.n890 AVDD.t574 1.60217
R2008 AVDD.n892 AVDD.t878 1.60217
R2009 AVDD.n894 AVDD.t303 1.60217
R2010 AVDD.n897 AVDD.t402 1.60217
R2011 AVDD.n899 AVDD.t386 1.60217
R2012 AVDD.n902 AVDD.t497 1.60217
R2013 AVDD.n892 AVDD.t978 1.60217
R2014 AVDD.n894 AVDD.t397 1.60217
R2015 AVDD.n897 AVDD.t513 1.60217
R2016 AVDD.n899 AVDD.t493 1.60217
R2017 AVDD.n902 AVDD.t614 1.60217
R2018 AVDD.n715 AVDD.t984 1.60217
R2019 AVDD.n743 AVDD.t181 1.60217
R2020 AVDD.n1179 AVDD.t724 1.60217
R2021 AVDD.n1006 AVDD.t1142 1.60217
R2022 AVDD.n1010 AVDD.t707 1.60217
R2023 AVDD.n982 AVDD.t817 1.60217
R2024 AVDD.n1096 AVDD.t246 1.60217
R2025 AVDD.n2101 AVDD.n2100 1.60175
R2026 AVDD.n1677 AVDD.n1676 1.60175
R2027 AVDD.n1214 AVDD.n1211 1.57603
R2028 AVDD.n1024 AVDD.n1021 1.57603
R2029 AVDD.n2109 AVDD.n46 1.5005
R2030 AVDD.n2074 AVDD.n2073 1.5005
R2031 AVDD.n2076 AVDD.n2075 1.5005
R2032 AVDD.n2133 AVDD.n2132 1.5005
R2033 AVDD.n2049 AVDD.n2048 1.5005
R2034 AVDD.n1854 AVDD.n1853 1.5005
R2035 AVDD.n1856 AVDD.n1855 1.5005
R2036 AVDD.n1922 AVDD.n1921 1.5005
R2037 AVDD.n1845 AVDD.n1844 1.5005
R2038 AVDD.n1887 AVDD.n67 1.5005
R2039 AVDD.n1641 AVDD.n1640 1.5005
R2040 AVDD.n1707 AVDD.n1706 1.5005
R2041 AVDD.n1662 AVDD.n1541 1.5005
R2042 AVDD.n1690 AVDD.n1689 1.5005
R2043 AVDD.n1709 AVDD.n1708 1.5005
R2044 AVDD.n263 AVDD.n185 1.5005
R2045 AVDD.n290 AVDD.n289 1.5005
R2046 AVDD.n341 AVDD.n340 1.5005
R2047 AVDD.n234 AVDD.n233 1.5005
R2048 AVDD.n339 AVDD.n338 1.5005
R2049 AVDD.n1726 AVDD.t1008 1.4705
R2050 AVDD.t138 AVDD.n1726 1.4705
R2051 AVDD.n162 AVDD.t1264 1.4705
R2052 AVDD.n162 AVDD.t1008 1.4705
R2053 AVDD.t422 AVDD.n166 1.4705
R2054 AVDD.n166 AVDD.t1264 1.4705
R2055 AVDD.n169 AVDD.t671 1.4705
R2056 AVDD.n169 AVDD.t384 1.4705
R2057 AVDD.t1076 AVDD.n174 1.4705
R2058 AVDD.n174 AVDD.t671 1.4705
R2059 AVDD.n177 AVDD.t111 1.4705
R2060 AVDD.n177 AVDD.t1108 1.4705
R2061 AVDD.t653 AVDD.n181 1.4705
R2062 AVDD.n181 AVDD.t111 1.4705
R2063 AVDD.n182 AVDD.t934 1.4705
R2064 AVDD.n182 AVDD.t653 1.4705
R2065 AVDD.n2137 AVDD.t948 1.4705
R2066 AVDD.t1208 AVDD.n2137 1.4705
R2067 AVDD.n1735 AVDD.t54 1.4705
R2068 AVDD.n1735 AVDD.t948 1.4705
R2069 AVDD.t1064 AVDD.n1739 1.4705
R2070 AVDD.n1739 AVDD.t54 1.4705
R2071 AVDD.n1742 AVDD.t713 1.4705
R2072 AVDD.n1742 AVDD.t1136 1.4705
R2073 AVDD.t418 AVDD.n1747 1.4705
R2074 AVDD.n1747 AVDD.t713 1.4705
R2075 AVDD.n1750 AVDD.t269 1.4705
R2076 AVDD.n1750 AVDD.t287 1.4705
R2077 AVDD.t643 AVDD.n1754 1.4705
R2078 AVDD.n1754 AVDD.t269 1.4705
R2079 AVDD.n1755 AVDD.t1168 1.4705
R2080 AVDD.n1755 AVDD.t643 1.4705
R2081 AVDD.t285 AVDD.n1319 1.4705
R2082 AVDD.n1319 AVDD.t665 1.4705
R2083 AVDD.n1320 AVDD.t966 1.4705
R2084 AVDD.n1320 AVDD.t285 1.4705
R2085 AVDD.t904 AVDD.n1324 1.4705
R2086 AVDD.n1324 AVDD.t966 1.4705
R2087 AVDD.n1327 AVDD.t906 1.4705
R2088 AVDD.n1327 AVDD.t527 1.4705
R2089 AVDD.t501 AVDD.n1332 1.4705
R2090 AVDD.n1332 AVDD.t906 1.4705
R2091 AVDD.t472 AVDD.n1337 1.4705
R2092 AVDD.n1337 AVDD.t90 1.4705
R2093 AVDD.n1338 AVDD.t748 1.4705
R2094 AVDD.n1338 AVDD.t472 1.4705
R2095 AVDD.t1098 AVDD.n1342 1.4705
R2096 AVDD.n1342 AVDD.t748 1.4705
R2097 AVDD.t1068 AVDD.n1355 1.4705
R2098 AVDD.n1355 AVDD.t1158 1.4705
R2099 AVDD.n1356 AVDD.t495 1.4705
R2100 AVDD.n1356 AVDD.t1068 1.4705
R2101 AVDD.t426 AVDD.n1360 1.4705
R2102 AVDD.n1360 AVDD.t495 1.4705
R2103 AVDD.n1363 AVDD.t98 1.4705
R2104 AVDD.n1363 AVDD.t1016 1.4705
R2105 AVDD.t6 AVDD.n1368 1.4705
R2106 AVDD.n1368 AVDD.t98 1.4705
R2107 AVDD.t1036 AVDD.n1373 1.4705
R2108 AVDD.n1373 AVDD.t594 1.4705
R2109 AVDD.n1374 AVDD.t1126 1.4705
R2110 AVDD.n1374 AVDD.t1036 1.4705
R2111 AVDD.t1210 AVDD.n1378 1.4705
R2112 AVDD.n1378 AVDD.t1126 1.4705
R2113 AVDD.n703 AVDD.t289 1.4705
R2114 AVDD.t673 AVDD.n703 1.4705
R2115 AVDD.n701 AVDD.t972 1.4705
R2116 AVDD.t289 AVDD.n701 1.4705
R2117 AVDD.n700 AVDD.t910 1.4705
R2118 AVDD.t972 AVDD.n700 1.4705
R2119 AVDD.n697 AVDD.t912 1.4705
R2120 AVDD.t533 AVDD.n697 1.4705
R2121 AVDD.n695 AVDD.t509 1.4705
R2122 AVDD.t912 AVDD.n695 1.4705
R2123 AVDD.n693 AVDD.t485 1.4705
R2124 AVDD.t102 AVDD.n693 1.4705
R2125 AVDD.n691 AVDD.t756 1.4705
R2126 AVDD.t485 AVDD.n691 1.4705
R2127 AVDD.n690 AVDD.t1104 1.4705
R2128 AVDD.t756 AVDD.n690 1.4705
R2129 AVDD.n685 AVDD.t1082 1.4705
R2130 AVDD.t1166 AVDD.n685 1.4705
R2131 AVDD.n683 AVDD.t503 1.4705
R2132 AVDD.t1082 AVDD.n683 1.4705
R2133 AVDD.n682 AVDD.t430 1.4705
R2134 AVDD.t503 AVDD.n682 1.4705
R2135 AVDD.n679 AVDD.t106 1.4705
R2136 AVDD.t1020 AVDD.n679 1.4705
R2137 AVDD.n678 AVDD.t11 1.4705
R2138 AVDD.t106 AVDD.n678 1.4705
R2139 AVDD.n676 AVDD.t1046 1.4705
R2140 AVDD.t600 AVDD.n676 1.4705
R2141 AVDD.n674 AVDD.t1134 1.4705
R2142 AVDD.t1046 AVDD.n674 1.4705
R2143 AVDD.n673 AVDD.t1216 1.4705
R2144 AVDD.t1134 AVDD.n673 1.4705
R2145 AVDD.n1287 AVDD.t766 1.4705
R2146 AVDD.t715 AVDD.n1287 1.4705
R2147 AVDD.n1282 AVDD.t1170 1.4705
R2148 AVDD.n1282 AVDD.t766 1.4705
R2149 AVDD.n1281 AVDD.t900 1.4705
R2150 AVDD.t1170 AVDD.n1281 1.4705
R2151 AVDD.n1276 AVDD.t186 1.4705
R2152 AVDD.t620 AVDD.n1276 1.4705
R2153 AVDD.n1271 AVDD.t239 1.4705
R2154 AVDD.n1271 AVDD.t186 1.4705
R2155 AVDD.n1268 AVDD.t37 1.4705
R2156 AVDD.t489 AVDD.n1268 1.4705
R2157 AVDD.n1263 AVDD.t628 1.4705
R2158 AVDD.n1263 AVDD.t37 1.4705
R2159 AVDD.n1262 AVDD.t206 1.4705
R2160 AVDD.t628 AVDD.n1262 1.4705
R2161 AVDD.n1948 AVDD.t869 1.4705
R2162 AVDD.t819 AVDD.n1948 1.4705
R2163 AVDD.n1944 AVDD.t1248 1.4705
R2164 AVDD.n1944 AVDD.t869 1.4705
R2165 AVDD.n1943 AVDD.t996 1.4705
R2166 AVDD.t1248 AVDD.n1943 1.4705
R2167 AVDD.n1938 AVDD.t305 1.4705
R2168 AVDD.t732 AVDD.n1938 1.4705
R2169 AVDD.n1933 AVDD.t343 1.4705
R2170 AVDD.n1933 AVDD.t305 1.4705
R2171 AVDD.n1930 AVDD.t145 1.4705
R2172 AVDD.t586 AVDD.n1930 1.4705
R2173 AVDD.n1926 AVDD.t738 1.4705
R2174 AVDD.n1926 AVDD.t145 1.4705
R2175 AVDD.n1925 AVDD.t311 1.4705
R2176 AVDD.t738 AVDD.n1925 1.4705
R2177 AVDD.n2043 AVDD.t1888 1.4705
R2178 AVDD.n2043 AVDD.n2042 1.4705
R2179 AVDD.n2045 AVDD.t1505 1.4705
R2180 AVDD.n2045 AVDD.n2044 1.4705
R2181 AVDD.n2005 AVDD.t1498 1.4705
R2182 AVDD.n2005 AVDD.n2004 1.4705
R2183 AVDD.n2007 AVDD.t1589 1.4705
R2184 AVDD.n2007 AVDD.n2006 1.4705
R2185 AVDD.n2121 AVDD.t1497 1.4705
R2186 AVDD.n2121 AVDD.n2120 1.4705
R2187 AVDD.n2124 AVDD.t1330 1.4705
R2188 AVDD.n2124 AVDD.n2123 1.4705
R2189 AVDD.n2127 AVDD.t1567 1.4705
R2190 AVDD.n2127 AVDD.n2126 1.4705
R2191 AVDD.n2130 AVDD.t1598 1.4705
R2192 AVDD.n2130 AVDD.n2129 1.4705
R2193 AVDD.n56 AVDD.t1514 1.4705
R2194 AVDD.n56 AVDD.n55 1.4705
R2195 AVDD.n53 AVDD.t1318 1.4705
R2196 AVDD.n53 AVDD.n52 1.4705
R2197 AVDD.n50 AVDD.t1614 1.4705
R2198 AVDD.n50 AVDD.n49 1.4705
R2199 AVDD.n48 AVDD.t1640 1.4705
R2200 AVDD.n48 AVDD.n47 1.4705
R2201 AVDD.n2097 AVDD.t1327 1.4705
R2202 AVDD.n2097 AVDD.n2096 1.4705
R2203 AVDD.n2091 AVDD.t1645 1.4705
R2204 AVDD.n2091 AVDD.n2090 1.4705
R2205 AVDD.n2085 AVDD.t1594 1.4705
R2206 AVDD.n2085 AVDD.n2084 1.4705
R2207 AVDD.n2079 AVDD.t1690 1.4705
R2208 AVDD.n2079 AVDD.n2078 1.4705
R2209 AVDD.n1976 AVDD.t1314 1.4705
R2210 AVDD.n1976 AVDD.n1975 1.4705
R2211 AVDD.n1970 AVDD.t1545 1.4705
R2212 AVDD.n1970 AVDD.n1969 1.4705
R2213 AVDD.n1964 AVDD.t1703 1.4705
R2214 AVDD.n1964 AVDD.n1963 1.4705
R2215 AVDD.n1961 AVDD.t1670 1.4705
R2216 AVDD.n1961 AVDD.n1960 1.4705
R2217 AVDD.n2062 AVDD.t1654 1.4705
R2218 AVDD.n2062 AVDD.n2061 1.4705
R2219 AVDD.n2065 AVDD.t1617 1.4705
R2220 AVDD.n2065 AVDD.n2064 1.4705
R2221 AVDD.n2068 AVDD.t1864 1.4705
R2222 AVDD.n2068 AVDD.n2067 1.4705
R2223 AVDD.n2071 AVDD.t1500 1.4705
R2224 AVDD.n2071 AVDD.n2070 1.4705
R2225 AVDD.n2059 AVDD.t1562 1.4705
R2226 AVDD.n2059 AVDD.n2058 1.4705
R2227 AVDD.n2056 AVDD.t1593 1.4705
R2228 AVDD.n2056 AVDD.n2055 1.4705
R2229 AVDD.n2053 AVDD.t1882 1.4705
R2230 AVDD.n2053 AVDD.n2052 1.4705
R2231 AVDD.n2051 AVDD.t1698 1.4705
R2232 AVDD.n2051 AVDD.n2050 1.4705
R2233 AVDD.n2035 AVDD.t1689 1.4705
R2234 AVDD.n2035 AVDD.n2034 1.4705
R2235 AVDD.n2029 AVDD.t1316 1.4705
R2236 AVDD.n2029 AVDD.n2028 1.4705
R2237 AVDD.n2023 AVDD.t1872 1.4705
R2238 AVDD.n2023 AVDD.n2022 1.4705
R2239 AVDD.n2017 AVDD.t1675 1.4705
R2240 AVDD.n2017 AVDD.n2016 1.4705
R2241 AVDD.n1999 AVDD.t1530 1.4705
R2242 AVDD.n1999 AVDD.n1998 1.4705
R2243 AVDD.n1993 AVDD.t1283 1.4705
R2244 AVDD.n1993 AVDD.n1992 1.4705
R2245 AVDD.n1987 AVDD.t1540 1.4705
R2246 AVDD.n1987 AVDD.n1986 1.4705
R2247 AVDD.n1984 AVDD.t1575 1.4705
R2248 AVDD.n1984 AVDD.n1983 1.4705
R2249 AVDD.n2111 AVDD.t1626 1.4705
R2250 AVDD.n2111 AVDD.n2110 1.4705
R2251 AVDD.n2113 AVDD.t1602 1.4705
R2252 AVDD.n2113 AVDD.n2112 1.4705
R2253 AVDD.n2103 AVDD.t1595 1.4705
R2254 AVDD.n2103 AVDD.n2102 1.4705
R2255 AVDD.n2105 AVDD.t1583 1.4705
R2256 AVDD.n2105 AVDD.n2104 1.4705
R2257 AVDD.n1778 AVDD.t1315 1.4705
R2258 AVDD.n1778 AVDD.n1777 1.4705
R2259 AVDD.n1788 AVDD.t1597 1.4705
R2260 AVDD.n1788 AVDD.n1787 1.4705
R2261 AVDD.n1865 AVDD.t1894 1.4705
R2262 AVDD.n1865 AVDD.n1864 1.4705
R2263 AVDD.n1867 AVDD.t1506 1.4705
R2264 AVDD.n1867 AVDD.n1866 1.4705
R2265 AVDD.n1870 AVDD.t1526 1.4705
R2266 AVDD.n1870 AVDD.n1869 1.4705
R2267 AVDD.n1872 AVDD.t1513 1.4705
R2268 AVDD.n1872 AVDD.n1871 1.4705
R2269 AVDD.n1876 AVDD.t1667 1.4705
R2270 AVDD.n1876 AVDD.n1875 1.4705
R2271 AVDD.n1878 AVDD.t1579 1.4705
R2272 AVDD.n1878 AVDD.n1877 1.4705
R2273 AVDD.n1882 AVDD.t1561 1.4705
R2274 AVDD.n1882 AVDD.n1881 1.4705
R2275 AVDD.n1884 AVDD.t1608 1.4705
R2276 AVDD.n1884 AVDD.n1883 1.4705
R2277 AVDD.n1889 AVDD.t1501 1.4705
R2278 AVDD.n1889 AVDD.n1888 1.4705
R2279 AVDD.n1891 AVDD.t1521 1.4705
R2280 AVDD.n1891 AVDD.n1890 1.4705
R2281 AVDD.n1895 AVDD.t1509 1.4705
R2282 AVDD.n1895 AVDD.n1894 1.4705
R2283 AVDD.n1897 AVDD.t1322 1.4705
R2284 AVDD.n1897 AVDD.n1896 1.4705
R2285 AVDD.n1901 AVDD.t1576 1.4705
R2286 AVDD.n1901 AVDD.n1900 1.4705
R2287 AVDD.n1903 AVDD.t1560 1.4705
R2288 AVDD.n1903 AVDD.n1902 1.4705
R2289 AVDD.n1907 AVDD.t1321 1.4705
R2290 AVDD.n1907 AVDD.n1906 1.4705
R2291 AVDD.n1909 AVDD.t1650 1.4705
R2292 AVDD.n1909 AVDD.n1908 1.4705
R2293 AVDD.n1822 AVDD.t1535 1.4705
R2294 AVDD.n1822 AVDD.n1821 1.4705
R2295 AVDD.n1824 AVDD.t1299 1.4705
R2296 AVDD.n1824 AVDD.n1823 1.4705
R2297 AVDD.n1827 AVDD.t1578 1.4705
R2298 AVDD.n1827 AVDD.n1826 1.4705
R2299 AVDD.n1829 AVDD.t1628 1.4705
R2300 AVDD.n1829 AVDD.n1828 1.4705
R2301 AVDD.n1833 AVDD.t1298 1.4705
R2302 AVDD.n1833 AVDD.n1832 1.4705
R2303 AVDD.n1835 AVDD.t1881 1.4705
R2304 AVDD.n1835 AVDD.n1834 1.4705
R2305 AVDD.n1839 AVDD.t1899 1.4705
R2306 AVDD.n1839 AVDD.n1838 1.4705
R2307 AVDD.n1841 AVDD.t1577 1.4705
R2308 AVDD.n1841 AVDD.n1840 1.4705
R2309 AVDD.n1816 AVDD.t1662 1.4705
R2310 AVDD.n1816 AVDD.n1815 1.4705
R2311 AVDD.n1818 AVDD.t1580 1.4705
R2312 AVDD.n1818 AVDD.n1817 1.4705
R2313 AVDD.n1810 AVDD.t1627 1.4705
R2314 AVDD.n1810 AVDD.n1809 1.4705
R2315 AVDD.n1812 AVDD.t1891 1.4705
R2316 AVDD.n1812 AVDD.n1811 1.4705
R2317 AVDD.n1804 AVDD.t1873 1.4705
R2318 AVDD.n1804 AVDD.n1803 1.4705
R2319 AVDD.n1806 AVDD.t1659 1.4705
R2320 AVDD.n1806 AVDD.n1805 1.4705
R2321 AVDD.n1798 AVDD.t1596 1.4705
R2322 AVDD.n1798 AVDD.n1797 1.4705
R2323 AVDD.n1800 AVDD.t1613 1.4705
R2324 AVDD.n1800 AVDD.n1799 1.4705
R2325 AVDD.n1919 AVDD.t1592 1.4705
R2326 AVDD.n1919 AVDD.n1918 1.4705
R2327 AVDD.n1915 AVDD.t1697 1.4705
R2328 AVDD.n1915 AVDD.n1914 1.4705
R2329 AVDD.n1770 AVDD.t1691 1.4705
R2330 AVDD.n1770 AVDD.n1769 1.4705
R2331 AVDD.n1764 AVDD.t1493 1.4705
R2332 AVDD.n1764 AVDD.n1763 1.4705
R2333 AVDD.n1851 AVDD.t1492 1.4705
R2334 AVDD.n1851 AVDD.n1850 1.4705
R2335 AVDD.n1847 AVDD.t1512 1.4705
R2336 AVDD.n1847 AVDD.n1846 1.4705
R2337 AVDD.t853 AVDD.n2167 1.4705
R2338 AVDD.n2167 AVDD.t1112 1.4705
R2339 AVDD.n2168 AVDD.t1242 1.4705
R2340 AVDD.n2168 AVDD.t853 1.4705
R2341 AVDD.t988 AVDD.n2172 1.4705
R2342 AVDD.n2172 AVDD.t1242 1.4705
R2343 AVDD.n2175 AVDD.t610 1.4705
R2344 AVDD.n2175 AVDD.t1024 1.4705
R2345 AVDD.t331 AVDD.n1387 1.4705
R2346 AVDD.n1387 AVDD.t610 1.4705
R2347 AVDD.t136 AVDD.n1392 1.4705
R2348 AVDD.n1392 AVDD.t153 1.4705
R2349 AVDD.n1393 AVDD.t549 1.4705
R2350 AVDD.n1393 AVDD.t136 1.4705
R2351 AVDD.t1056 AVDD.n1397 1.4705
R2352 AVDD.n1397 AVDD.t549 1.4705
R2353 AVDD.n31 AVDD.t188 1.4705
R2354 AVDD.t466 AVDD.n31 1.4705
R2355 AVDD.n29 AVDD.t618 1.4705
R2356 AVDD.t188 AVDD.n29 1.4705
R2357 AVDD.n28 AVDD.t341 1.4705
R2358 AVDD.t618 AVDD.n28 1.4705
R2359 AVDD.t1228 AVDD.n25 1.4705
R2360 AVDD.t376 AVDD.n25 1.4705
R2361 AVDD.t964 AVDD.n1385 1.4705
R2362 AVDD.n1385 AVDD.t1228 1.4705
R2363 AVDD.n1384 AVDD.t800 1.4705
R2364 AVDD.t813 AVDD.n1384 1.4705
R2365 AVDD.n1382 AVDD.t1174 1.4705
R2366 AVDD.t800 AVDD.n1382 1.4705
R2367 AVDD.n1381 AVDD.t412 1.4705
R2368 AVDD.t1174 AVDD.n1381 1.4705
R2369 AVDD.n552 AVDD.t1164 1.4705
R2370 AVDD.t736 AVDD.n552 1.4705
R2371 AVDD.n547 AVDD.t280 1.4705
R2372 AVDD.n547 AVDD.t1164 1.4705
R2373 AVDD.n546 AVDD.t699 1.4705
R2374 AVDD.t280 AVDD.n546 1.4705
R2375 AVDD.n541 AVDD.t1234 1.4705
R2376 AVDD.t970 AVDD.n541 1.4705
R2377 AVDD.n536 AVDD.t382 1.4705
R2378 AVDD.n536 AVDD.t1234 1.4705
R2379 AVDD.n533 AVDD.t624 1.4705
R2380 AVDD.t348 AVDD.n533 1.4705
R2381 AVDD.n528 AVDD.t940 1.4705
R2382 AVDD.n528 AVDD.t624 1.4705
R2383 AVDD.n527 AVDD.t1200 1.4705
R2384 AVDD.t940 AVDD.n527 1.4705
R2385 AVDD.n550 AVDD.t292 1.4705
R2386 AVDD.n550 AVDD.t1140 1.4705
R2387 AVDD.n549 AVDD.t675 1.4705
R2388 AVDD.t292 AVDD.n549 1.4705
R2389 AVDD.n544 AVDD.t1078 1.4705
R2390 AVDD.n544 AVDD.t675 1.4705
R2391 AVDD.n539 AVDD.t364 1.4705
R2392 AVDD.n539 AVDD.t60 1.4705
R2393 AVDD.n538 AVDD.t804 1.4705
R2394 AVDD.t364 AVDD.n538 1.4705
R2395 AVDD.n531 AVDD.t1022 1.4705
R2396 AVDD.n531 AVDD.t758 1.4705
R2397 AVDD.n530 AVDD.t20 1.4705
R2398 AVDD.t1022 AVDD.n530 1.4705
R2399 AVDD.n525 AVDD.t333 1.4705
R2400 AVDD.n525 AVDD.t20 1.4705
R2401 AVDD.t119 AVDD.n465 1.4705
R2402 AVDD.n465 AVDD.t558 1.4705
R2403 AVDD.n466 AVDD.t400 1.4705
R2404 AVDD.n466 AVDD.t119 1.4705
R2405 AVDD.t839 AVDD.n470 1.4705
R2406 AVDD.n470 AVDD.t400 1.4705
R2407 AVDD.n473 AVDD.t1052 1.4705
R2408 AVDD.n473 AVDD.t796 1.4705
R2409 AVDD.t201 AVDD.n478 1.4705
R2410 AVDD.n478 AVDD.t1052 1.4705
R2411 AVDD.t505 AVDD.n483 1.4705
R2412 AVDD.n483 AVDD.t227 1.4705
R2413 AVDD.n484 AVDD.t1030 1.4705
R2414 AVDD.n484 AVDD.t505 1.4705
R2415 AVDD.t1280 AVDD.n488 1.4705
R2416 AVDD.n488 AVDD.t1030 1.4705
R2417 AVDD.n462 AVDD.t523 1.4705
R2418 AVDD.n462 AVDD.t950 1.4705
R2419 AVDD.n460 AVDD.t815 1.4705
R2420 AVDD.t523 AVDD.n460 1.4705
R2421 AVDD.n459 AVDD.t1218 1.4705
R2422 AVDD.t815 AVDD.n459 1.4705
R2423 AVDD.n456 AVDD.t175 1.4705
R2424 AVDD.t1176 AVDD.n456 1.4705
R2425 AVDD.n455 AVDD.t612 1.4705
R2426 AVDD.t175 AVDD.n455 1.4705
R2427 AVDD.n453 AVDD.t916 1.4705
R2428 AVDD.t630 AVDD.n453 1.4705
R2429 AVDD.n451 AVDD.t148 1.4705
R2430 AVDD.t916 AVDD.n451 1.4705
R2431 AVDD.n450 AVDD.t434 1.4705
R2432 AVDD.t148 AVDD.n450 1.4705
R2433 AVDD.t1040 AVDD.n1468 1.4705
R2434 AVDD.n1468 AVDD.t454 1.4705
R2435 AVDD.n1469 AVDD.t1110 1.4705
R2436 AVDD.n1469 AVDD.t1040 1.4705
R2437 AVDD.t762 AVDD.n1473 1.4705
R2438 AVDD.n1473 AVDD.t1110 1.4705
R2439 AVDD.n1476 AVDD.t231 1.4705
R2440 AVDD.n1476 AVDD.t156 1.4705
R2441 AVDD.n666 AVDD.t1146 1.4705
R2442 AVDD.t231 AVDD.n666 1.4705
R2443 AVDD.n661 AVDD.t535 1.4705
R2444 AVDD.t462 AVDD.n661 1.4705
R2445 AVDD.n656 AVDD.t164 1.4705
R2446 AVDD.n656 AVDD.t535 1.4705
R2447 AVDD.n655 AVDD.t244 1.4705
R2448 AVDD.t164 AVDD.n655 1.4705
R2449 AVDD.n645 AVDD.t786 1.4705
R2450 AVDD.t1148 AVDD.n645 1.4705
R2451 AVDD.n640 AVDD.t857 1.4705
R2452 AVDD.n640 AVDD.t786 1.4705
R2453 AVDD.n639 AVDD.t460 1.4705
R2454 AVDD.t857 AVDD.n639 1.4705
R2455 AVDD.n634 AVDD.t908 1.4705
R2456 AVDD.t859 AVDD.n634 1.4705
R2457 AVDD.n629 AVDD.t531 1.4705
R2458 AVDD.n629 AVDD.t908 1.4705
R2459 AVDD.n626 AVDD.t1270 1.4705
R2460 AVDD.t1224 AVDD.n626 1.4705
R2461 AVDD.n621 AVDD.t768 1.4705
R2462 AVDD.n621 AVDD.t1270 1.4705
R2463 AVDD.n620 AVDD.t821 1.4705
R2464 AVDD.t768 AVDD.n620 1.4705
R2465 AVDD.n671 AVDD.t1048 1.4705
R2466 AVDD.t464 AVDD.n671 1.4705
R2467 AVDD.n669 AVDD.t1118 1.4705
R2468 AVDD.t1048 AVDD.n669 1.4705
R2469 AVDD.n668 AVDD.t770 1.4705
R2470 AVDD.t1118 AVDD.n668 1.4705
R2471 AVDD.t236 AVDD.n123 1.4705
R2472 AVDD.t160 AVDD.n123 1.4705
R2473 AVDD.t1152 AVDD.n663 1.4705
R2474 AVDD.n663 AVDD.t236 1.4705
R2475 AVDD.n659 AVDD.t541 1.4705
R2476 AVDD.n659 AVDD.t474 1.4705
R2477 AVDD.n658 AVDD.t172 1.4705
R2478 AVDD.t541 AVDD.n658 1.4705
R2479 AVDD.n653 AVDD.t250 1.4705
R2480 AVDD.n653 AVDD.t172 1.4705
R2481 AVDD.n643 AVDD.t788 1.4705
R2482 AVDD.n643 AVDD.t1156 1.4705
R2483 AVDD.n642 AVDD.t865 1.4705
R2484 AVDD.t788 AVDD.n642 1.4705
R2485 AVDD.n637 AVDD.t468 1.4705
R2486 AVDD.n637 AVDD.t865 1.4705
R2487 AVDD.n632 AVDD.t914 1.4705
R2488 AVDD.n632 AVDD.t861 1.4705
R2489 AVDD.n631 AVDD.t539 1.4705
R2490 AVDD.t914 AVDD.n631 1.4705
R2491 AVDD.n624 AVDD.t1274 1.4705
R2492 AVDD.n624 AVDD.t1230 1.4705
R2493 AVDD.n623 AVDD.t772 1.4705
R2494 AVDD.t1274 AVDD.n623 1.4705
R2495 AVDD.n618 AVDD.t829 1.4705
R2496 AVDD.n618 AVDD.t772 1.4705
R2497 AVDD.t689 AVDD.n573 1.4705
R2498 AVDD.n573 AVDD.t275 1.4705
R2499 AVDD.n574 AVDD.t1062 1.4705
R2500 AVDD.n574 AVDD.t689 1.4705
R2501 AVDD.t218 AVDD.n578 1.4705
R2502 AVDD.n578 AVDD.t1062 1.4705
R2503 AVDD.n581 AVDD.t792 1.4705
R2504 AVDD.n581 AVDD.t491 1.4705
R2505 AVDD.t1190 AVDD.n586 1.4705
R2506 AVDD.n586 AVDD.t792 1.4705
R2507 AVDD.t133 AVDD.n591 1.4705
R2508 AVDD.n591 AVDD.t1160 1.4705
R2509 AVDD.n592 AVDD.t446 1.4705
R2510 AVDD.n592 AVDD.t133 1.4705
R2511 AVDD.t750 AVDD.n596 1.4705
R2512 AVDD.n596 AVDD.t446 1.4705
R2513 AVDD.t944 AVDD.n424 1.4705
R2514 AVDD.n424 AVDD.t51 1.4705
R2515 AVDD.n425 AVDD.t1202 1.4705
R2516 AVDD.n425 AVDD.t944 1.4705
R2517 AVDD.t360 AVDD.n429 1.4705
R2518 AVDD.n429 AVDD.t1202 1.4705
R2519 AVDD.n432 AVDD.t590 1.4705
R2520 AVDD.n432 AVDD.t317 1.4705
R2521 AVDD.t1012 AVDD.n437 1.4705
R2522 AVDD.n437 AVDD.t590 1.4705
R2523 AVDD.t1278 AVDD.n442 1.4705
R2524 AVDD.n442 AVDD.t1028 1.4705
R2525 AVDD.n443 AVDD.t580 1.4705
R2526 AVDD.n443 AVDD.t1278 1.4705
R2527 AVDD.t873 AVDD.n447 1.4705
R2528 AVDD.n447 AVDD.t580 1.4705
R2529 AVDD.t661 AVDD.n1509 1.4705
R2530 AVDD.n1509 AVDD.t242 1.4705
R2531 AVDD.n1510 AVDD.t1034 1.4705
R2532 AVDD.n1510 AVDD.t661 1.4705
R2533 AVDD.t193 AVDD.n1514 1.4705
R2534 AVDD.n1514 AVDD.t1034 1.4705
R2535 AVDD.n1517 AVDD.t764 1.4705
R2536 AVDD.n1517 AVDD.t456 1.4705
R2537 AVDD.t1172 AVDD.n382 1.4705
R2538 AVDD.n382 AVDD.t764 1.4705
R2539 AVDD.t122 AVDD.n387 1.4705
R2540 AVDD.n387 AVDD.t1128 1.4705
R2541 AVDD.n388 AVDD.t424 1.4705
R2542 AVDD.n388 AVDD.t122 1.4705
R2543 AVDD.t728 AVDD.n392 1.4705
R2544 AVDD.n392 AVDD.t424 1.4705
R2545 AVDD.n108 AVDD.t1268 1.4705
R2546 AVDD.t886 AVDD.n108 1.4705
R2547 AVDD.n106 AVDD.t404 1.4705
R2548 AVDD.t1268 AVDD.n106 1.4705
R2549 AVDD.n105 AVDD.t847 1.4705
R2550 AVDD.t404 AVDD.n105 1.4705
R2551 AVDD.t88 AVDD.n102 1.4705
R2552 AVDD.t1092 AVDD.n102 1.4705
R2553 AVDD.t525 AVDD.n380 1.4705
R2554 AVDD.n380 AVDD.t88 1.4705
R2555 AVDD.n379 AVDD.t778 1.4705
R2556 AVDD.t483 AVDD.n379 1.4705
R2557 AVDD.n377 AVDD.t1058 1.4705
R2558 AVDD.t778 AVDD.n377 1.4705
R2559 AVDD.n376 AVDD.t45 1.4705
R2560 AVDD.t1058 AVDD.n376 1.4705
R2561 AVDD.n1537 AVDD.t780 1.4705
R2562 AVDD.t345 AVDD.n1537 1.4705
R2563 AVDD.n1533 AVDD.t1162 1.4705
R2564 AVDD.n1533 AVDD.t780 1.4705
R2565 AVDD.n1532 AVDD.t307 1.4705
R2566 AVDD.t1162 AVDD.n1532 1.4705
R2567 AVDD.n1527 AVDD.t871 1.4705
R2568 AVDD.t576 AVDD.n1527 1.4705
R2569 AVDD.t1254 AVDD.n350 1.4705
R2570 AVDD.n350 AVDD.t871 1.4705
R2571 AVDD.t224 AVDD.n355 1.4705
R2572 AVDD.n355 AVDD.t1214 1.4705
R2573 AVDD.n356 AVDD.t537 1.4705
R2574 AVDD.n356 AVDD.t224 1.4705
R2575 AVDD.t827 AVDD.n360 1.4705
R2576 AVDD.n360 AVDD.t537 1.4705
R2577 AVDD.n1643 AVDD.t1843 1.4705
R2578 AVDD.n1643 AVDD.n1642 1.4705
R2579 AVDD.n1645 AVDD.t1437 1.4705
R2580 AVDD.n1645 AVDD.n1644 1.4705
R2581 AVDD.n1583 AVDD.t1808 1.4705
R2582 AVDD.n1583 AVDD.n1582 1.4705
R2583 AVDD.n1585 AVDD.t1406 1.4705
R2584 AVDD.n1585 AVDD.n1584 1.4705
R2585 AVDD.n1720 AVDD.t1381 1.4705
R2586 AVDD.n1720 AVDD.n1719 1.4705
R2587 AVDD.n1717 AVDD.t1793 1.4705
R2588 AVDD.n1717 AVDD.n1716 1.4705
R2589 AVDD.n1714 AVDD.t1450 1.4705
R2590 AVDD.n1714 AVDD.n1713 1.4705
R2591 AVDD.n1711 AVDD.t1395 1.4705
R2592 AVDD.n1711 AVDD.n1710 1.4705
R2593 AVDD.n83 AVDD.t1422 1.4705
R2594 AVDD.n83 AVDD.n82 1.4705
R2595 AVDD.n80 AVDD.t1832 1.4705
R2596 AVDD.n80 AVDD.n79 1.4705
R2597 AVDD.n77 AVDD.t1844 1.4705
R2598 AVDD.n77 AVDD.n76 1.4705
R2599 AVDD.n75 AVDD.t1412 1.4705
R2600 AVDD.n75 AVDD.n74 1.4705
R2601 AVDD.n1579 AVDD.t1342 1.4705
R2602 AVDD.n1579 AVDD.n1578 1.4705
R2603 AVDD.n1575 AVDD.t1761 1.4705
R2604 AVDD.n1575 AVDD.n1574 1.4705
R2605 AVDD.n1571 AVDD.t1835 1.4705
R2606 AVDD.n1571 AVDD.n1570 1.4705
R2607 AVDD.n1567 AVDD.t1358 1.4705
R2608 AVDD.n1567 AVDD.n1566 1.4705
R2609 AVDD.n1561 AVDD.t1396 1.4705
R2610 AVDD.n1561 AVDD.n1560 1.4705
R2611 AVDD.n1555 AVDD.t1790 1.4705
R2612 AVDD.n1555 AVDD.n1554 1.4705
R2613 AVDD.n1549 AVDD.t1812 1.4705
R2614 AVDD.n1549 AVDD.n1548 1.4705
R2615 AVDD.n1546 AVDD.t1386 1.4705
R2616 AVDD.n1546 AVDD.n1545 1.4705
R2617 AVDD.n1673 AVDD.t1839 1.4705
R2618 AVDD.n1673 AVDD.n1672 1.4705
R2619 AVDD.n1670 AVDD.t1389 1.4705
R2620 AVDD.n1670 AVDD.n1669 1.4705
R2621 AVDD.n1667 AVDD.t1756 1.4705
R2622 AVDD.n1667 AVDD.n1666 1.4705
R2623 AVDD.n1664 AVDD.t1850 1.4705
R2624 AVDD.n1664 AVDD.n1663 1.4705
R2625 AVDD.n1660 AVDD.t1469 1.4705
R2626 AVDD.n1660 AVDD.n1659 1.4705
R2627 AVDD.n1657 AVDD.t1407 1.4705
R2628 AVDD.n1657 AVDD.n1656 1.4705
R2629 AVDD.n1654 AVDD.t1423 1.4705
R2630 AVDD.n1654 AVDD.n1653 1.4705
R2631 AVDD.n1652 AVDD.t1458 1.4705
R2632 AVDD.n1652 AVDD.n1651 1.4705
R2633 AVDD.n1626 AVDD.t1480 1.4705
R2634 AVDD.n1626 AVDD.n1625 1.4705
R2635 AVDD.n1622 AVDD.t1394 1.4705
R2636 AVDD.n1622 AVDD.n1621 1.4705
R2637 AVDD.n1618 AVDD.t1428 1.4705
R2638 AVDD.n1618 AVDD.n1617 1.4705
R2639 AVDD.n1614 AVDD.t1792 1.4705
R2640 AVDD.n1614 AVDD.n1613 1.4705
R2641 AVDD.n1608 AVDD.t1388 1.4705
R2642 AVDD.n1608 AVDD.n1607 1.4705
R2643 AVDD.n1602 AVDD.t1747 1.4705
R2644 AVDD.n1602 AVDD.n1601 1.4705
R2645 AVDD.n1596 AVDD.t1847 1.4705
R2646 AVDD.n1596 AVDD.n1595 1.4705
R2647 AVDD.n1593 AVDD.t1380 1.4705
R2648 AVDD.n1593 AVDD.n1592 1.4705
R2649 AVDD.n1701 AVDD.t1385 1.4705
R2650 AVDD.n1701 AVDD.n1700 1.4705
R2651 AVDD.n1703 AVDD.t1371 1.4705
R2652 AVDD.n1703 AVDD.n1702 1.4705
R2653 AVDD.n1692 AVDD.t1343 1.4705
R2654 AVDD.n1692 AVDD.n1691 1.4705
R2655 AVDD.n1694 AVDD.t1483 1.4705
R2656 AVDD.n1694 AVDD.n1693 1.4705
R2657 AVDD.n228 AVDD.t1805 1.4705
R2658 AVDD.n228 AVDD.n227 1.4705
R2659 AVDD.n220 AVDD.t1356 1.4705
R2660 AVDD.n220 AVDD.n219 1.4705
R2661 AVDD.n316 AVDD.t1398 1.4705
R2662 AVDD.n316 AVDD.n315 1.4705
R2663 AVDD.n318 AVDD.t1387 1.4705
R2664 AVDD.n318 AVDD.n317 1.4705
R2665 AVDD.n321 AVDD.t1827 1.4705
R2666 AVDD.n321 AVDD.n320 1.4705
R2667 AVDD.n323 AVDD.t1811 1.4705
R2668 AVDD.n323 AVDD.n322 1.4705
R2669 AVDD.n327 AVDD.t1472 1.4705
R2670 AVDD.n327 AVDD.n326 1.4705
R2671 AVDD.n329 AVDD.t1456 1.4705
R2672 AVDD.n329 AVDD.n328 1.4705
R2673 AVDD.n333 AVDD.t1409 1.4705
R2674 AVDD.n333 AVDD.n332 1.4705
R2675 AVDD.n335 AVDD.t1399 1.4705
R2676 AVDD.n335 AVDD.n334 1.4705
R2677 AVDD.n310 AVDD.t1754 1.4705
R2678 AVDD.n310 AVDD.n309 1.4705
R2679 AVDD.n312 AVDD.t1433 1.4705
R2680 AVDD.n312 AVDD.n311 1.4705
R2681 AVDD.n304 AVDD.t1849 1.4705
R2682 AVDD.n304 AVDD.n303 1.4705
R2683 AVDD.n306 AVDD.t1840 1.4705
R2684 AVDD.n306 AVDD.n305 1.4705
R2685 AVDD.n298 AVDD.t1449 1.4705
R2686 AVDD.n298 AVDD.n297 1.4705
R2687 AVDD.n300 AVDD.t1848 1.4705
R2688 AVDD.n300 AVDD.n299 1.4705
R2689 AVDD.n292 AVDD.t1740 1.4705
R2690 AVDD.n292 AVDD.n291 1.4705
R2691 AVDD.n294 AVDD.t1418 1.4705
R2692 AVDD.n294 AVDD.n293 1.4705
R2693 AVDD.n190 AVDD.t1444 1.4705
R2694 AVDD.n190 AVDD.n189 1.4705
R2695 AVDD.n192 AVDD.t1455 1.4705
R2696 AVDD.n192 AVDD.n191 1.4705
R2697 AVDD.n195 AVDD.t1402 1.4705
R2698 AVDD.n195 AVDD.n194 1.4705
R2699 AVDD.n197 AVDD.t1372 1.4705
R2700 AVDD.n197 AVDD.n196 1.4705
R2701 AVDD.n201 AVDD.t1779 1.4705
R2702 AVDD.n201 AVDD.n200 1.4705
R2703 AVDD.n203 AVDD.t1405 1.4705
R2704 AVDD.n203 AVDD.n202 1.4705
R2705 AVDD.n207 AVDD.t1457 1.4705
R2706 AVDD.n207 AVDD.n206 1.4705
R2707 AVDD.n209 AVDD.t1769 1.4705
R2708 AVDD.n209 AVDD.n208 1.4705
R2709 AVDD.n236 AVDD.t1339 1.4705
R2710 AVDD.n236 AVDD.n235 1.4705
R2711 AVDD.n238 AVDD.t1364 1.4705
R2712 AVDD.n238 AVDD.n237 1.4705
R2713 AVDD.n242 AVDD.t1434 1.4705
R2714 AVDD.n242 AVDD.n241 1.4705
R2715 AVDD.n244 AVDD.t1419 1.4705
R2716 AVDD.n244 AVDD.n243 1.4705
R2717 AVDD.n248 AVDD.t1755 1.4705
R2718 AVDD.n248 AVDD.n247 1.4705
R2719 AVDD.n250 AVDD.t1826 1.4705
R2720 AVDD.n250 AVDD.n249 1.4705
R2721 AVDD.n254 AVDD.t1484 1.4705
R2722 AVDD.n254 AVDD.n253 1.4705
R2723 AVDD.n256 AVDD.t1349 1.4705
R2724 AVDD.n256 AVDD.n255 1.4705
R2725 AVDD.n153 AVDD.t1359 1.4705
R2726 AVDD.n153 AVDD.n152 1.4705
R2727 AVDD.n344 AVDD.t1475 1.4705
R2728 AVDD.n344 AVDD.n343 1.4705
R2729 AVDD.n285 AVDD.t1408 1.4705
R2730 AVDD.n285 AVDD.n284 1.4705
R2731 AVDD.n277 AVDD.t1379 1.4705
R2732 AVDD.n277 AVDD.n276 1.4705
R2733 AVDD.n261 AVDD.t1823 1.4705
R2734 AVDD.n261 AVDD.n260 1.4705
R2735 AVDD.n266 AVDD.t1780 1.4705
R2736 AVDD.n266 AVDD.n265 1.4705
R2737 AVDD.n1437 AVDD.t918 1.4705
R2738 AVDD.t23 AVDD.n1437 1.4705
R2739 AVDD.n1432 AVDD.t1182 1.4705
R2740 AVDD.n1432 AVDD.t918 1.4705
R2741 AVDD.n1431 AVDD.t339 1.4705
R2742 AVDD.t1182 AVDD.n1431 1.4705
R2743 AVDD.n1426 AVDD.t568 1.4705
R2744 AVDD.t299 AVDD.n1426 1.4705
R2745 AVDD.n1421 AVDD.t994 1.4705
R2746 AVDD.n1421 AVDD.t568 1.4705
R2747 AVDD.n1418 AVDD.t1266 1.4705
R2748 AVDD.t1010 AVDD.n1418 1.4705
R2749 AVDD.n1413 AVDD.t560 1.4705
R2750 AVDD.n1413 AVDD.t1266 1.4705
R2751 AVDD.n1412 AVDD.t845 1.4705
R2752 AVDD.t560 AVDD.n1412 1.4705
R2753 AVDD.n1435 AVDD.t277 1.4705
R2754 AVDD.n1435 AVDD.t693 1.4705
R2755 AVDD.n1434 AVDD.t553 1.4705
R2756 AVDD.t277 AVDD.n1434 1.4705
R2757 AVDD.n1429 AVDD.t974 1.4705
R2758 AVDD.n1429 AVDD.t553 1.4705
R2759 AVDD.n1424 AVDD.t1194 1.4705
R2760 AVDD.n1424 AVDD.t928 1.4705
R2761 AVDD.n1423 AVDD.t352 1.4705
R2762 AVDD.t1194 AVDD.n1423 1.4705
R2763 AVDD.n1416 AVDD.t649 1.4705
R2764 AVDD.n1416 AVDD.t369 1.4705
R2765 AVDD.n1415 AVDD.t1180 1.4705
R2766 AVDD.t649 AVDD.n1415 1.4705
R2767 AVDD.n1410 AVDD.t178 1.4705
R2768 AVDD.n1410 AVDD.t1180 1.4705
R2769 AVDD.n1228 AVDD.t1186 1.4705
R2770 AVDD.n1228 AVDD.t790 1.4705
R2771 AVDD.n1227 AVDD.t922 1.4705
R2772 AVDD.t1186 AVDD.n1227 1.4705
R2773 AVDD.t216 AVDD.n776 1.4705
R2774 AVDD.n776 AVDD.t641 1.4705
R2775 AVDD.n777 AVDD.t273 1.4705
R2776 AVDD.n777 AVDD.t216 1.4705
R2777 AVDD.t65 AVDD.n949 1.4705
R2778 AVDD.n949 AVDD.t511 1.4705
R2779 AVDD.n950 AVDD.t657 1.4705
R2780 AVDD.n950 AVDD.t65 1.4705
R2781 AVDD.n940 AVDD.t229 1.4705
R2782 AVDD.n940 AVDD.t657 1.4705
R2783 AVDD.n923 AVDD.t880 1.4705
R2784 AVDD.t1154 AVDD.n923 1.4705
R2785 AVDD.n771 AVDD.t744 1.4705
R2786 AVDD.n771 AVDD.t1204 1.4705
R2787 AVDD.n766 AVDD.t367 1.4705
R2788 AVDD.t744 AVDD.n766 1.4705
R2789 AVDD.t1252 AVDD.n780 1.4705
R2790 AVDD.n780 AVDD.t367 1.4705
R2791 AVDD.n944 AVDD.t1122 1.4705
R2792 AVDD.t1044 AVDD.n944 1.4705
R2793 AVDD.n943 AVDD.t28 1.4705
R2794 AVDD.t1122 AVDD.n943 1.4705
R2795 AVDD.n937 AVDD.t902 1.4705
R2796 AVDD.t687 AVDD.n937 1.4705
R2797 AVDD.n931 AVDD.t962 1.4705
R2798 AVDD.n931 AVDD.t902 1.4705
R2799 AVDD.n930 AVDD.t476 1.4705
R2800 AVDD.t962 AVDD.n930 1.4705
R2801 AVDD.n1232 AVDD.t790 1.4705
R2802 AVDD.t740 AVDD.n1232 1.4705
R2803 AVDD.n919 AVDD.t1260 1.4705
R2804 AVDD.t880 AVDD.n919 1.4705
R2805 AVDD.n913 AVDD.t1006 1.4705
R2806 AVDD.n913 AVDD.t1260 1.4705
R2807 AVDD.n910 AVDD.t632 1.4705
R2808 AVDD.t1042 AVDD.n910 1.4705
R2809 AVDD.t356 AVDD.n2184 1.4705
R2810 AVDD.n2184 AVDD.t632 1.4705
R2811 AVDD.t170 AVDD.n2189 1.4705
R2812 AVDD.n2189 AVDD.t183 1.4705
R2813 AVDD.n2190 AVDD.t572 1.4705
R2814 AVDD.n2190 AVDD.t170 1.4705
R2815 AVDD.t1074 AVDD.n2194 1.4705
R2816 AVDD.n2194 AVDD.t572 1.4705
R2817 AVDD.n878 AVDD.t31 1.4705
R2818 AVDD.t336 AVDD.n878 1.4705
R2819 AVDD.n873 AVDD.t470 1.4705
R2820 AVDD.n873 AVDD.t31 1.4705
R2821 AVDD.n872 AVDD.t196 1.4705
R2822 AVDD.t470 AVDD.n872 1.4705
R2823 AVDD.n867 AVDD.t1086 1.4705
R2824 AVDD.t253 AVDD.n867 1.4705
R2825 AVDD.n862 AVDD.t835 1.4705
R2826 AVDD.n862 AVDD.t1086 1.4705
R2827 AVDD.n859 AVDD.t645 1.4705
R2828 AVDD.t663 AVDD.n859 1.4705
R2829 AVDD.n854 AVDD.t1026 1.4705
R2830 AVDD.n854 AVDD.t645 1.4705
R2831 AVDD.n853 AVDD.t295 1.4705
R2832 AVDD.t1026 AVDD.n853 1.4705
R2833 AVDD.n876 AVDD.t444 1.4705
R2834 AVDD.n876 AVDD.t746 1.4705
R2835 AVDD.n875 AVDD.t892 1.4705
R2836 AVDD.t444 AVDD.n875 1.4705
R2837 AVDD.n870 AVDD.t602 1.4705
R2838 AVDD.n870 AVDD.t892 1.4705
R2839 AVDD.n865 AVDD.t220 1.4705
R2840 AVDD.n865 AVDD.t647 1.4705
R2841 AVDD.n864 AVDD.t1212 1.4705
R2842 AVDD.t220 AVDD.n864 1.4705
R2843 AVDD.n857 AVDD.t1032 1.4705
R2844 AVDD.n857 AVDD.t1054 1.4705
R2845 AVDD.n856 AVDD.t141 1.4705
R2846 AVDD.t1032 AVDD.n856 1.4705
R2847 AVDD.n851 AVDD.t683 1.4705
R2848 AVDD.n851 AVDD.t141 1.4705
R2849 AVDD.t1232 AVDD.n814 1.4705
R2850 AVDD.n814 AVDD.t1198 1.4705
R2851 AVDD.n815 AVDD.t379 1.4705
R2852 AVDD.n815 AVDD.t1232 1.4705
R2853 AVDD.t93 AVDD.n819 1.4705
R2854 AVDD.n819 AVDD.t379 1.4705
R2855 AVDD.n822 AVDD.t697 1.4705
R2856 AVDD.n822 AVDD.t1102 1.4705
R2857 AVDD.t734 AVDD.n827 1.4705
R2858 AVDD.n827 AVDD.t697 1.4705
R2859 AVDD.t562 AVDD.n832 1.4705
R2860 AVDD.n832 AVDD.t986 1.4705
R2861 AVDD.n833 AVDD.t1124 1.4705
R2862 AVDD.n833 AVDD.t562 1.4705
R2863 AVDD.t709 AVDD.n837 1.4705
R2864 AVDD.n837 AVDD.t1124 1.4705
R2865 AVDD.n800 AVDD.t362 1.4705
R2866 AVDD.t326 AVDD.n800 1.4705
R2867 AVDD.n798 AVDD.t802 1.4705
R2868 AVDD.t362 AVDD.n798 1.4705
R2869 AVDD.n797 AVDD.t507 1.4705
R2870 AVDD.t802 AVDD.n797 1.4705
R2871 AVDD.n794 AVDD.t1072 1.4705
R2872 AVDD.t234 AVDD.n794 1.4705
R2873 AVDD.n793 AVDD.t1138 1.4705
R2874 AVDD.t1072 AVDD.n793 1.4705
R2875 AVDD.n791 AVDD.t956 1.4705
R2876 AVDD.t83 AVDD.n791 1.4705
R2877 AVDD.n789 AVDD.t256 1.4705
R2878 AVDD.t956 AVDD.n789 1.4705
R2879 AVDD.n788 AVDD.t1088 1.4705
R2880 AVDD.t256 AVDD.n788 1.4705
R2881 AVDD.n1220 AVDD.t1720 1.4705
R2882 AVDD.n1220 AVDD.n1219 1.4705
R2883 AVDD.n1217 AVDD.t1704 1.4705
R2884 AVDD.n1217 AVDD.n1216 1.4705
R2885 AVDD.n1213 AVDD.t1646 1.4705
R2886 AVDD.n1213 AVDD.n1212 1.4705
R2887 AVDD.n1210 AVDD.t1726 1.4705
R2888 AVDD.n1210 AVDD.n1209 1.4705
R2889 AVDD.n1207 AVDD.t1713 1.4705
R2890 AVDD.n1207 AVDD.n1206 1.4705
R2891 AVDD.n739 AVDD.t1325 1.4705
R2892 AVDD.n739 AVDD.n738 1.4705
R2893 AVDD.n735 AVDD.t1601 1.4705
R2894 AVDD.n735 AVDD.n734 1.4705
R2895 AVDD.n731 AVDD.t1574 1.4705
R2896 AVDD.n731 AVDD.n730 1.4705
R2897 AVDD.n724 AVDD.t1629 1.4705
R2898 AVDD.n724 AVDD.n723 1.4705
R2899 AVDD.n720 AVDD.t1880 1.4705
R2900 AVDD.n720 AVDD.n719 1.4705
R2901 AVDD.n1172 AVDD.t1605 1.4705
R2902 AVDD.n1172 AVDD.n1171 1.4705
R2903 AVDD.n1175 AVDD.t1853 1.4705
R2904 AVDD.n1175 AVDD.n1174 1.4705
R2905 AVDD.n1164 AVDD.t1504 1.4705
R2906 AVDD.n1164 AVDD.n1163 1.4705
R2907 AVDD.n1167 AVDD.t1544 1.4705
R2908 AVDD.n1167 AVDD.n1166 1.4705
R2909 AVDD.n1156 AVDD.t1725 1.4705
R2910 AVDD.n1156 AVDD.n1155 1.4705
R2911 AVDD.n1159 AVDD.t1705 1.4705
R2912 AVDD.n1159 AVDD.n1158 1.4705
R2913 AVDD.n1142 AVDD.t1693 1.4705
R2914 AVDD.n1142 AVDD.n1141 1.4705
R2915 AVDD.n1145 AVDD.t1494 1.4705
R2916 AVDD.n1145 AVDD.n1144 1.4705
R2917 AVDD.n1134 AVDD.t1674 1.4705
R2918 AVDD.n1134 AVDD.n1133 1.4705
R2919 AVDD.n1137 AVDD.t1692 1.4705
R2920 AVDD.n1137 AVDD.n1136 1.4705
R2921 AVDD.n1013 AVDD.t1606 1.4705
R2922 AVDD.n1013 AVDD.n1012 1.4705
R2923 AVDD.n1016 AVDD.t1729 1.4705
R2924 AVDD.n1016 AVDD.n1015 1.4705
R2925 AVDD.n1020 AVDD.t1491 1.4705
R2926 AVDD.n1020 AVDD.n1019 1.4705
R2927 AVDD.n1023 AVDD.t1694 1.4705
R2928 AVDD.n1023 AVDD.n1022 1.4705
R2929 AVDD.n1026 AVDD.t1676 1.4705
R2930 AVDD.n1026 AVDD.n1025 1.4705
R2931 AVDD.n980 AVDD.t1716 1.4705
R2932 AVDD.n980 AVDD.n979 1.4705
R2933 AVDD.n976 AVDD.t1798 1.4705
R2934 AVDD.n976 AVDD.n975 1.4705
R2935 AVDD.n972 AVDD.t1885 1.4705
R2936 AVDD.n972 AVDD.n971 1.4705
R2937 AVDD.n965 AVDD.t1719 1.4705
R2938 AVDD.n965 AVDD.n964 1.4705
R2939 AVDD.n961 AVDD.t1710 1.4705
R2940 AVDD.n961 AVDD.n960 1.4705
R2941 AVDD.n1094 AVDD.t324 1.4705
R2942 AVDD.t811 AVDD.n1094 1.4705
R2943 AVDD.n1090 AVDD.t1222 1.4705
R2944 AVDD.n1090 AVDD.t324 1.4705
R2945 AVDD.n1089 AVDD.t876 1.4705
R2946 AVDD.t1222 AVDD.n1089 1.4705
R2947 AVDD.n1084 AVDD.t718 1.4705
R2948 AVDD.t639 AVDD.n1084 1.4705
R2949 AVDD.n1079 AVDD.t926 1.4705
R2950 AVDD.n1079 AVDD.t718 1.4705
R2951 AVDD.n1076 AVDD.t481 1.4705
R2952 AVDD.t283 AVDD.n1076 1.4705
R2953 AVDD.n1072 AVDD.t556 1.4705
R2954 AVDD.n1072 AVDD.t481 1.4705
R2955 AVDD.n1071 AVDD.t40 1.4705
R2956 AVDD.t556 AVDD.n1071 1.4705
R2957 AVDD.n1285 AVDD.t85 1.4705
R2958 AVDD.n1285 AVDD.t34 1.4705
R2959 AVDD.n1284 AVDD.t519 1.4705
R2960 AVDD.t85 AVDD.n1284 1.4705
R2961 AVDD.n1279 AVDD.t258 1.4705
R2962 AVDD.n1279 AVDD.t519 1.4705
R2963 AVDD.n1274 AVDD.t841 1.4705
R2964 AVDD.n1274 AVDD.t1240 1.4705
R2965 AVDD.n1273 AVDD.t884 1.4705
R2966 AVDD.t841 AVDD.n1273 1.4705
R2967 AVDD.n1266 AVDD.t705 1.4705
R2968 AVDD.n1266 AVDD.t1114 1.4705
R2969 AVDD.n1265 AVDD.t1244 1.4705
R2970 AVDD.t705 AVDD.n1265 1.4705
R2971 AVDD.n1260 AVDD.t851 1.4705
R2972 AVDD.n1260 AVDD.t1244 1.4705
R2973 AVDD.n2041 AVDD.n2040 1.46537
R2974 AVDD.n2047 AVDD.n2046 1.46537
R2975 AVDD.n2010 AVDD.n2009 1.46537
R2976 AVDD.n2117 AVDD.n2116 1.46537
R2977 AVDD.n2115 AVDD.n2114 1.46537
R2978 AVDD.n2108 AVDD.n2107 1.46537
R2979 AVDD.n1649 AVDD.n1648 1.46537
R2980 AVDD.n1647 AVDD.n1646 1.46537
R2981 AVDD.n1588 AVDD.n1587 1.46537
R2982 AVDD.n1699 AVDD.n1698 1.46537
R2983 AVDD.n1705 AVDD.n1704 1.46537
R2984 AVDD.n1697 AVDD.n1696 1.46537
R2985 AVDD.n1874 AVDD.n1873 1.46537
R2986 AVDD.n1880 AVDD.n1879 1.46537
R2987 AVDD.n1886 AVDD.n1885 1.46537
R2988 AVDD.n1893 AVDD.n1892 1.46537
R2989 AVDD.n1899 AVDD.n1898 1.46537
R2990 AVDD.n1905 AVDD.n1904 1.46537
R2991 AVDD.n1911 AVDD.n1910 1.46537
R2992 AVDD.n1831 AVDD.n1830 1.46537
R2993 AVDD.n1837 AVDD.n1836 1.46537
R2994 AVDD.n1843 AVDD.n1842 1.46537
R2995 AVDD.n1820 AVDD.n1819 1.46537
R2996 AVDD.n1814 AVDD.n1813 1.46537
R2997 AVDD.n1808 AVDD.n1807 1.46537
R2998 AVDD.n1802 AVDD.n1801 1.46537
R2999 AVDD.n325 AVDD.n324 1.46537
R3000 AVDD.n331 AVDD.n330 1.46537
R3001 AVDD.n337 AVDD.n336 1.46537
R3002 AVDD.n314 AVDD.n313 1.46537
R3003 AVDD.n308 AVDD.n307 1.46537
R3004 AVDD.n302 AVDD.n301 1.46537
R3005 AVDD.n296 AVDD.n295 1.46537
R3006 AVDD.n199 AVDD.n198 1.46537
R3007 AVDD.n205 AVDD.n204 1.46537
R3008 AVDD.n211 AVDD.n210 1.46537
R3009 AVDD.n240 AVDD.n239 1.46537
R3010 AVDD.n246 AVDD.n245 1.46537
R3011 AVDD.n252 AVDD.n251 1.46537
R3012 AVDD.n258 AVDD.n257 1.46537
R3013 AVDD.n1188 AVDD.n1187 1.30325
R3014 AVDD.n1162 AVDD.n1161 1.30325
R3015 AVDD.n1105 AVDD.n1104 1.30325
R3016 AVDD.n1221 AVDD.n1218 1.27338
R3017 AVDD.n1211 AVDD.n1208 1.27338
R3018 AVDD.n1215 AVDD.n1214 1.27228
R3019 AVDD.n1027 AVDD.n1024 1.27228
R3020 AVDD.n1021 AVDD.n1018 1.27228
R3021 AVDD.n1017 AVDD.n1014 1.27228
R3022 AVDD.n57 AVDD.n54 1.27228
R3023 AVDD.n2131 AVDD.n2128 1.27228
R3024 AVDD.n2125 AVDD.n2122 1.27228
R3025 AVDD.n2060 AVDD.n2057 1.27228
R3026 AVDD.n2072 AVDD.n2069 1.27228
R3027 AVDD.n2066 AVDD.n2063 1.27228
R3028 AVDD.n2117 AVDD.n2115 1.27228
R3029 AVDD.n2047 AVDD.n2041 1.27228
R3030 AVDD.n1911 AVDD.n1905 1.27228
R3031 AVDD.n1899 AVDD.n1893 1.27228
R3032 AVDD.n1886 AVDD.n1880 1.27228
R3033 AVDD.n1808 AVDD.n1802 1.27228
R3034 AVDD.n1820 AVDD.n1814 1.27228
R3035 AVDD.n1843 AVDD.n1837 1.27228
R3036 AVDD.n1917 AVDD.n1916 1.27228
R3037 AVDD.n1849 AVDD.n1848 1.27228
R3038 AVDD.n84 AVDD.n81 1.27228
R3039 AVDD.n1715 AVDD.n1712 1.27228
R3040 AVDD.n1721 AVDD.n1718 1.27228
R3041 AVDD.n1661 AVDD.n1658 1.27228
R3042 AVDD.n1668 AVDD.n1665 1.27228
R3043 AVDD.n1674 AVDD.n1671 1.27228
R3044 AVDD.n1705 AVDD.n1699 1.27228
R3045 AVDD.n1649 AVDD.n1647 1.27228
R3046 AVDD.n302 AVDD.n296 1.27228
R3047 AVDD.n314 AVDD.n308 1.27228
R3048 AVDD.n337 AVDD.n331 1.27228
R3049 AVDD.n258 AVDD.n252 1.27228
R3050 AVDD.n246 AVDD.n240 1.27228
R3051 AVDD.n211 AVDD.n205 1.27228
R3052 AVDD.n345 AVDD.n342 1.27228
R3053 AVDD.n267 AVDD.n264 1.27228
R3054 AVDD.n1522 AVDD.t87 1.1382
R3055 AVDD.n1481 AVDD.t174 1.1382
R3056 AVDD.n2180 AVDD.t97 1.1382
R3057 AVDD.n1126 AVDD.t185 1.1382
R3058 AVDD.n2135 AVDD.n2134 1.13692
R3059 AVDD.n1951 AVDD.n58 1.13692
R3060 AVDD.n1724 AVDD.n1723 1.13692
R3061 AVDD.n1540 AVDD.n85 1.13692
R3062 AVDD.n1974 AVDD.n1973 0.9995
R3063 AVDD.n2083 AVDD.n2082 0.9995
R3064 AVDD.n2095 AVDD.n2094 0.9995
R3065 AVDD.n1997 AVDD.n1996 0.9995
R3066 AVDD.n2021 AVDD.n2020 0.9995
R3067 AVDD.n2033 AVDD.n2032 0.9995
R3068 AVDD.n1559 AVDD.n1558 0.9995
R3069 AVDD.n1686 AVDD.n1685 0.9995
R3070 AVDD.n1680 AVDD.n1679 0.9995
R3071 AVDD.n1606 AVDD.n1605 0.9995
R3072 AVDD.n1636 AVDD.n1635 0.9995
R3073 AVDD.n1630 AVDD.n1629 0.9995
R3074 AVDD.n1197 AVDD.n1196 0.9995
R3075 AVDD.n1191 AVDD.n1190 0.9995
R3076 AVDD.n1185 AVDD.n1184 0.9995
R3077 AVDD.n1140 AVDD.n1139 0.9995
R3078 AVDD.n1154 AVDD.n1153 0.9995
R3079 AVDD.n1170 AVDD.n1169 0.9995
R3080 AVDD.n1114 AVDD.n1113 0.9995
R3081 AVDD.n1108 AVDD.n1107 0.9995
R3082 AVDD.n1102 AVDD.n1101 0.9995
R3083 AVDD.n1860 AVDD.n1859 0.991625
R3084 AVDD.n1793 AVDD.n1792 0.991625
R3085 AVDD.n275 AVDD.n274 0.991625
R3086 AVDD.n218 AVDD.n217 0.991625
R3087 AVDD.n2134 AVDD.n2133 0.983405
R3088 AVDD.n2119 AVDD.n1951 0.983405
R3089 AVDD.n1723 AVDD.n1722 0.983405
R3090 AVDD.n1708 AVDD.n1540 0.983405
R3091 AVDD.n1218 AVDD.n1215 0.937025
R3092 AVDD.n1018 AVDD.n1017 0.937025
R3093 AVDD.n2075 AVDD.n2074 0.822966
R3094 AVDD.n2101 AVDD.n1952 0.822966
R3095 AVDD.n1676 AVDD.n1675 0.822966
R3096 AVDD.n1690 AVDD.n1541 0.822966
R3097 AVDD.n1913 AVDD.n1912 0.737223
R3098 AVDD.n1796 AVDD.n1758 0.737223
R3099 AVDD.n1922 AVDD.n67 0.737223
R3100 AVDD.n1854 AVDD.n1845 0.737223
R3101 AVDD.n340 AVDD.n339 0.737223
R3102 AVDD.n233 AVDD.n185 0.737223
R3103 AVDD.n346 AVDD.n151 0.737223
R3104 AVDD.n268 AVDD.n259 0.737223
R3105 AVDD.n1863 AVDD.n1758 0.725061
R3106 AVDD.n1855 AVDD.n1854 0.725061
R3107 AVDD.n290 AVDD.n185 0.725061
R3108 AVDD.n269 AVDD.n268 0.725061
R3109 AVDD.n1194 AVDD.n1193 0.66425
R3110 AVDD.n1148 AVDD.n1147 0.66425
R3111 AVDD.n1111 AVDD.n1110 0.66425
R3112 AVDD.n2133 AVDD.n46 0.639318
R3113 AVDD.n2074 AVDD.n2049 0.639318
R3114 AVDD.n2119 AVDD.n2118 0.639318
R3115 AVDD.n2039 AVDD.n1952 0.639318
R3116 AVDD.n1722 AVDD.n73 0.639318
R3117 AVDD.n1675 AVDD.n1650 0.639318
R3118 AVDD.n1708 AVDD.n1707 0.639318
R3119 AVDD.n1640 AVDD.n1541 0.639318
R3120 AVDD.n2075 AVDD.n46 0.585196
R3121 AVDD.n2118 AVDD.n2101 0.585196
R3122 AVDD.n1912 AVDD.n1863 0.585196
R3123 AVDD.n1855 AVDD.n67 0.585196
R3124 AVDD.n1676 AVDD.n73 0.585196
R3125 AVDD.n1707 AVDD.n1690 0.585196
R3126 AVDD.n339 AVDD.n290 0.585196
R3127 AVDD.n269 AVDD.n151 0.585196
R3128 AVDD.n2132 AVDD.n57 0.236091
R3129 AVDD.n2073 AVDD.n2060 0.236091
R3130 AVDD.n1709 AVDD.n84 0.236091
R3131 AVDD.n1662 AVDD.n1661 0.236091
R3132 AVDD.n1050 AVDD.n1049 0.166289
R3133 AVDD.n1122 AVDD.n1121 0.166289
R3134 AVDD.n1123 AVDD.n1122 0.166289
R3135 AVDD.n1887 AVDD.n1886 0.150184
R3136 AVDD.n1844 AVDD.n1843 0.150184
R3137 AVDD.n338 AVDD.n337 0.150184
R3138 AVDD.n234 AVDD.n211 0.150184
R3139 AVDD.n1962 AVDD.n1959 0.14
R3140 AVDD.n1967 AVDD.n1959 0.14
R3141 AVDD.n1968 AVDD.n1958 0.14
R3142 AVDD.n1973 AVDD.n1958 0.14
R3143 AVDD.n1974 AVDD.n1957 0.14
R3144 AVDD.n1979 AVDD.n1957 0.14
R3145 AVDD.n2077 AVDD.n1956 0.14
R3146 AVDD.n2082 AVDD.n1956 0.14
R3147 AVDD.n2083 AVDD.n1955 0.14
R3148 AVDD.n2088 AVDD.n1955 0.14
R3149 AVDD.n2089 AVDD.n1954 0.14
R3150 AVDD.n2094 AVDD.n1954 0.14
R3151 AVDD.n2095 AVDD.n1953 0.14
R3152 AVDD.n2100 AVDD.n1953 0.14
R3153 AVDD.n1985 AVDD.n1982 0.14
R3154 AVDD.n1990 AVDD.n1982 0.14
R3155 AVDD.n1991 AVDD.n1981 0.14
R3156 AVDD.n1996 AVDD.n1981 0.14
R3157 AVDD.n1997 AVDD.n1980 0.14
R3158 AVDD.n2002 AVDD.n1980 0.14
R3159 AVDD.n2015 AVDD.n2014 0.14
R3160 AVDD.n2020 AVDD.n2014 0.14
R3161 AVDD.n2021 AVDD.n2013 0.14
R3162 AVDD.n2026 AVDD.n2013 0.14
R3163 AVDD.n2027 AVDD.n2012 0.14
R3164 AVDD.n2032 AVDD.n2012 0.14
R3165 AVDD.n2033 AVDD.n2011 0.14
R3166 AVDD.n2038 AVDD.n2011 0.14
R3167 AVDD.n1862 AVDD.n1759 0.14
R3168 AVDD.n1860 AVDD.n1759 0.14
R3169 AVDD.n1859 AVDD.n1762 0.14
R3170 AVDD.n1857 AVDD.n1762 0.14
R3171 AVDD.n1773 AVDD.n1766 0.14
R3172 AVDD.n1771 AVDD.n1766 0.14
R3173 AVDD.n1795 AVDD.n1783 0.14
R3174 AVDD.n1793 AVDD.n1783 0.14
R3175 AVDD.n1792 AVDD.n1786 0.14
R3176 AVDD.n1790 AVDD.n1786 0.14
R3177 AVDD.n1781 AVDD.n1774 0.14
R3178 AVDD.n1779 AVDD.n1774 0.14
R3179 AVDD.n1547 AVDD.n1544 0.14
R3180 AVDD.n1552 AVDD.n1544 0.14
R3181 AVDD.n1553 AVDD.n1543 0.14
R3182 AVDD.n1558 AVDD.n1543 0.14
R3183 AVDD.n1559 AVDD.n1542 0.14
R3184 AVDD.n1564 AVDD.n1542 0.14
R3185 AVDD.n1688 AVDD.n1565 0.14
R3186 AVDD.n1686 AVDD.n1565 0.14
R3187 AVDD.n1685 AVDD.n1569 0.14
R3188 AVDD.n1683 AVDD.n1569 0.14
R3189 AVDD.n1682 AVDD.n1573 0.14
R3190 AVDD.n1680 AVDD.n1573 0.14
R3191 AVDD.n1679 AVDD.n1577 0.14
R3192 AVDD.n1677 AVDD.n1577 0.14
R3193 AVDD.n1594 AVDD.n1591 0.14
R3194 AVDD.n1599 AVDD.n1591 0.14
R3195 AVDD.n1600 AVDD.n1590 0.14
R3196 AVDD.n1605 AVDD.n1590 0.14
R3197 AVDD.n1606 AVDD.n1589 0.14
R3198 AVDD.n1611 AVDD.n1589 0.14
R3199 AVDD.n1638 AVDD.n1612 0.14
R3200 AVDD.n1636 AVDD.n1612 0.14
R3201 AVDD.n1635 AVDD.n1616 0.14
R3202 AVDD.n1633 AVDD.n1616 0.14
R3203 AVDD.n1632 AVDD.n1620 0.14
R3204 AVDD.n1630 AVDD.n1620 0.14
R3205 AVDD.n1629 AVDD.n1624 0.14
R3206 AVDD.n1624 AVDD.n1581 0.14
R3207 AVDD.n270 AVDD.n187 0.14
R3208 AVDD.n274 AVDD.n187 0.14
R3209 AVDD.n275 AVDD.n186 0.14
R3210 AVDD.n280 AVDD.n186 0.14
R3211 AVDD.n288 AVDD.n281 0.14
R3212 AVDD.n286 AVDD.n281 0.14
R3213 AVDD.n213 AVDD.n188 0.14
R3214 AVDD.n217 AVDD.n213 0.14
R3215 AVDD.n218 AVDD.n212 0.14
R3216 AVDD.n223 AVDD.n212 0.14
R3217 AVDD.n231 AVDD.n224 0.14
R3218 AVDD.n229 AVDD.n224 0.14
R3219 AVDD.n1199 AVDD.n718 0.14
R3220 AVDD.n1197 AVDD.n718 0.14
R3221 AVDD.n1196 AVDD.n722 0.14
R3222 AVDD.n1194 AVDD.n722 0.14
R3223 AVDD.n1193 AVDD.n726 0.14
R3224 AVDD.n1191 AVDD.n726 0.14
R3225 AVDD.n1190 AVDD.n729 0.14
R3226 AVDD.n1188 AVDD.n729 0.14
R3227 AVDD.n1187 AVDD.n733 0.14
R3228 AVDD.n1185 AVDD.n733 0.14
R3229 AVDD.n1184 AVDD.n737 0.14
R3230 AVDD.n1182 AVDD.n737 0.14
R3231 AVDD.n1132 AVDD.n750 0.14
R3232 AVDD.n1139 AVDD.n750 0.14
R3233 AVDD.n1140 AVDD.n749 0.14
R3234 AVDD.n1147 AVDD.n749 0.14
R3235 AVDD.n1148 AVDD.n748 0.14
R3236 AVDD.n1153 AVDD.n748 0.14
R3237 AVDD.n1154 AVDD.n747 0.14
R3238 AVDD.n1161 AVDD.n747 0.14
R3239 AVDD.n1162 AVDD.n746 0.14
R3240 AVDD.n1169 AVDD.n746 0.14
R3241 AVDD.n1170 AVDD.n745 0.14
R3242 AVDD.n1177 AVDD.n745 0.14
R3243 AVDD.n1116 AVDD.n959 0.14
R3244 AVDD.n1114 AVDD.n959 0.14
R3245 AVDD.n1113 AVDD.n963 0.14
R3246 AVDD.n1111 AVDD.n963 0.14
R3247 AVDD.n1110 AVDD.n967 0.14
R3248 AVDD.n1108 AVDD.n967 0.14
R3249 AVDD.n1107 AVDD.n970 0.14
R3250 AVDD.n1105 AVDD.n970 0.14
R3251 AVDD.n1104 AVDD.n974 0.14
R3252 AVDD.n1102 AVDD.n974 0.14
R3253 AVDD.n1101 AVDD.n978 0.14
R3254 AVDD.n1099 AVDD.n978 0.14
R3255 AVDD.n998 AVDD.n955 0.13175
R3256 AVDD.n1048 AVDD.n955 0.13175
R3257 AVDD.n994 AVDD.n956 0.13175
R3258 AVDD.n1048 AVDD.n956 0.13175
R3259 AVDD.n1243 AVDD.n1242 0.105779
R3260 AVDD.n1236 AVDD.n1235 0.105779
R3261 AVDD.n364 AVDD.n363 0.103153
R3262 AVDD.n600 AVDD.n599 0.103153
R3263 AVDD.n1300 AVDD.n1299 0.101802
R3264 AVDD.n808 AVDD.n804 0.101802
R3265 AVDD.n1299 AVDD.n1298 0.101802
R3266 AVDD.n1313 AVDD.n705 0.101802
R3267 AVDD.n1313 AVDD.n1312 0.101802
R3268 AVDD.n808 AVDD.n807 0.101802
R3269 AVDD.n2076 AVDD.n1979 0.10175
R3270 AVDD.n2003 AVDD.n2002 0.10175
R3271 AVDD.n1689 AVDD.n1564 0.10175
R3272 AVDD.n1639 AVDD.n1611 0.10175
R3273 AVDD.n396 AVDD.n373 0.0992755
R3274 AVDD.n397 AVDD.n396 0.0992755
R3275 AVDD.n614 AVDD.n406 0.0992755
R3276 AVDD.n614 AVDD.n613 0.0992755
R3277 AVDD.n521 AVDD.n517 0.0992755
R3278 AVDD.n521 AVDD.n520 0.0992755
R3279 AVDD.n606 AVDD.n605 0.0931471
R3280 AVDD.n607 AVDD.n606 0.0931471
R3281 AVDD.n562 AVDD.n561 0.0931471
R3282 AVDD.n561 AVDD.n114 0.0931471
R3283 AVDD.n562 AVDD.n115 0.0931471
R3284 AVDD.n1496 AVDD.n115 0.0931471
R3285 AVDD.n898 AVDD.n20 0.0931471
R3286 AVDD.n37 AVDD.n20 0.0931471
R3287 AVDD.n898 AVDD.n38 0.0931471
R3288 AVDD.n2154 AVDD.n38 0.0931471
R3289 AVDD.n1241 AVDD.n1240 0.0931471
R3290 AVDD.n1306 AVDD.n1241 0.0931471
R3291 AVDD.n609 AVDD.n608 0.0931471
R3292 AVDD.n608 AVDD.n607 0.0931471
R3293 AVDD.n494 AVDD.n493 0.0931471
R3294 AVDD.n493 AVDD.n114 0.0931471
R3295 AVDD.n494 AVDD.n116 0.0931471
R3296 AVDD.n1496 AVDD.n116 0.0931471
R3297 AVDD.n884 AVDD.n883 0.0931471
R3298 AVDD.n883 AVDD.n37 0.0931471
R3299 AVDD.n884 AVDD.n39 0.0931471
R3300 AVDD.n2154 AVDD.n39 0.0931471
R3301 AVDD.n401 AVDD.n99 0.0931471
R3302 AVDD.n607 AVDD.n99 0.0931471
R3303 AVDD.n1498 AVDD.n100 0.0931471
R3304 AVDD.n114 AVDD.n100 0.0931471
R3305 AVDD.n1498 AVDD.n1497 0.0931471
R3306 AVDD.n1497 AVDD.n1496 0.0931471
R3307 AVDD.n369 AVDD.n91 0.0931471
R3308 AVDD.n607 AVDD.n91 0.0931471
R3309 AVDD.n1494 AVDD.n92 0.0931471
R3310 AVDD.n114 AVDD.n92 0.0931471
R3311 AVDD.n1495 AVDD.n1494 0.0931471
R3312 AVDD.n1496 AVDD.n1495 0.0931471
R3313 AVDD.n1305 AVDD.n1304 0.0931471
R3314 AVDD.n1306 AVDD.n1305 0.0931471
R3315 AVDD.n1294 AVDD.n708 0.0931471
R3316 AVDD.n1306 AVDD.n708 0.0931471
R3317 AVDD.n1308 AVDD.n1307 0.0931471
R3318 AVDD.n1307 AVDD.n1306 0.0931471
R3319 AVDD.n2156 AVDD.n23 0.0931471
R3320 AVDD.n37 AVDD.n23 0.0931471
R3321 AVDD.n2156 AVDD.n2155 0.0931471
R3322 AVDD.n2155 AVDD.n2154 0.0931471
R3323 AVDD.n2152 AVDD.n2146 0.0931471
R3324 AVDD.n2146 AVDD.n37 0.0931471
R3325 AVDD.n2153 AVDD.n2152 0.0931471
R3326 AVDD.n2154 AVDD.n2153 0.0931471
R3327 AVDD.n2203 AVDD.n14 0.0931471
R3328 AVDD.n14 AVDD.n5 0.0931471
R3329 AVDD.n2203 AVDD.n7 0.0931471
R3330 AVDD.n2219 AVDD.n7 0.0931471
R3331 AVDD.n2217 AVDD.n11 0.0931471
R3332 AVDD.n11 AVDD.n5 0.0931471
R3333 AVDD.n2218 AVDD.n2217 0.0931471
R3334 AVDD.n2219 AVDD.n2218 0.0931471
R3335 AVDD.n1452 AVDD.n1451 0.0931471
R3336 AVDD.n1451 AVDD.n5 0.0931471
R3337 AVDD.n1452 AVDD.n6 0.0931471
R3338 AVDD.n2219 AVDD.n6 0.0931471
R3339 AVDD.n2221 AVDD.n1 0.0931471
R3340 AVDD.n5 AVDD.n1 0.0931471
R3341 AVDD.n2221 AVDD.n2220 0.0931471
R3342 AVDD.n2220 AVDD.n2219 0.0931471
R3343 AVDD.n1130 AVDD.n1129 0.0737558
R3344 AVDD.n1129 AVDD.n1128 0.0737558
R3345 AVDD.n1124 AVDD.n744 0.0737558
R3346 AVDD.n1304 AVDD.n1303 0.0723953
R3347 AVDD.n1240 AVDD.n1239 0.0723953
R3348 AVDD.n1294 AVDD.n1293 0.0723953
R3349 AVDD.n1308 AVDD.n706 0.0723953
R3350 AVDD.n1059 AVDD.n1057 0.0720299
R3351 AVDD.n370 AVDD.n369 0.070602
R3352 AVDD.n1098 AVDD.n1097 0.0692176
R3353 AVDD.n953 AVDD.n952 0.0682419
R3354 AVDD.n1125 AVDD.n953 0.0682419
R3355 AVDD.n1081 AVDD.n954 0.0682419
R3356 AVDD.n1125 AVDD.n954 0.0682419
R3357 AVDD.n508 AVDD.n97 0.0682419
R3358 AVDD.n1522 AVDD.n97 0.0682419
R3359 AVDD.n476 AVDD.n121 0.0682419
R3360 AVDD.n1481 AVDD.n121 0.0682419
R3361 AVDD.n846 AVDD.n22 0.0682419
R3362 AVDD.n2180 AVDD.n22 0.0682419
R3363 AVDD.n825 AVDD.n709 0.0682419
R3364 AVDD.n1126 AVDD.n709 0.0682419
R3365 AVDD.n142 AVDD.n98 0.0682419
R3366 AVDD.n1522 AVDD.n98 0.0682419
R3367 AVDD.n1480 AVDD.n1479 0.0682419
R3368 AVDD.n1481 AVDD.n1480 0.0682419
R3369 AVDD.n1521 AVDD.n1520 0.0682419
R3370 AVDD.n1522 AVDD.n1521 0.0682419
R3371 AVDD.n118 AVDD.n112 0.0682419
R3372 AVDD.n1481 AVDD.n112 0.0682419
R3373 AVDD.n2179 AVDD.n2178 0.0682419
R3374 AVDD.n2180 AVDD.n2179 0.0682419
R3375 AVDD.n1524 AVDD.n1523 0.0682419
R3376 AVDD.n1523 AVDD.n1522 0.0682419
R3377 AVDD.n1935 AVDD.n40 0.0682419
R3378 AVDD.n1126 AVDD.n40 0.0682419
R3379 AVDD.n1255 AVDD.n35 0.0682419
R3380 AVDD.n1126 AVDD.n35 0.0682419
R3381 AVDD.n1366 AVDD.n8 0.0682419
R3382 AVDD.n2180 AVDD.n8 0.0682419
R3383 AVDD.n1330 AVDD.n696 0.0682419
R3384 AVDD.n1126 AVDD.n696 0.0682419
R3385 AVDD.n1745 AVDD.n3 0.0682419
R3386 AVDD.n2180 AVDD.n3 0.0682419
R3387 AVDD.n172 AVDD.n117 0.0682419
R3388 AVDD.n1481 AVDD.n117 0.0682419
R3389 AVDD.n584 AVDD.n96 0.0668158
R3390 AVDD.n1522 AVDD.n96 0.0668158
R3391 AVDD.n435 AVDD.n120 0.0668158
R3392 AVDD.n1481 AVDD.n120 0.0668158
R3393 AVDD.n2182 AVDD.n2181 0.0668158
R3394 AVDD.n2181 AVDD.n2180 0.0668158
R3395 AVDD.n762 AVDD.n710 0.0668158
R3396 AVDD.n1126 AVDD.n710 0.0668158
R3397 AVDD.n508 AVDD.n95 0.0668158
R3398 AVDD.n1522 AVDD.n95 0.0668158
R3399 AVDD.n476 AVDD.n119 0.0668158
R3400 AVDD.n1481 AVDD.n119 0.0668158
R3401 AVDD.n846 AVDD.n9 0.0668158
R3402 AVDD.n2180 AVDD.n9 0.0668158
R3403 AVDD.n825 AVDD.n707 0.0668158
R3404 AVDD.n1126 AVDD.n707 0.0668158
R3405 AVDD.n142 AVDD.n94 0.0668158
R3406 AVDD.n1522 AVDD.n94 0.0668158
R3407 AVDD.n1479 AVDD.n113 0.0668158
R3408 AVDD.n1481 AVDD.n113 0.0668158
R3409 AVDD.n1520 AVDD.n93 0.0668158
R3410 AVDD.n1522 AVDD.n93 0.0668158
R3411 AVDD.n1482 AVDD.n118 0.0668158
R3412 AVDD.n1482 AVDD.n1481 0.0668158
R3413 AVDD.n2178 AVDD.n4 0.0668158
R3414 AVDD.n2180 AVDD.n4 0.0668158
R3415 AVDD.n1255 AVDD.n41 0.0668158
R3416 AVDD.n1126 AVDD.n41 0.0668158
R3417 AVDD.n1366 AVDD.n21 0.0668158
R3418 AVDD.n2180 AVDD.n21 0.0668158
R3419 AVDD.n1330 AVDD.n36 0.0668158
R3420 AVDD.n1126 AVDD.n36 0.0668158
R3421 AVDD.n403 AVDD.n402 0.0660102
R3422 AVDD.n514 AVDD.n407 0.0660102
R3423 AVDD.n1304 AVDD.n1246 0.0629767
R3424 AVDD.n1240 AVDD.n711 0.0629767
R3425 AVDD.n1295 AVDD.n1294 0.0629767
R3426 AVDD.n1309 AVDD.n1308 0.0629767
R3427 AVDD.n1224 AVDD.n1222 0.0619118
R3428 AVDD.n1205 AVDD.n716 0.0616241
R3429 AVDD.n401 AVDD.n400 0.0614184
R3430 AVDD.n610 AVDD.n609 0.0614184
R3431 AVDD.n605 AVDD.n408 0.0614184
R3432 AVDD.n1485 AVDD.n1484 0.0525345
R3433 AVDD.n1490 AVDD.n1489 0.0525345
R3434 AVDD.n1503 AVDD.n1502 0.0525345
R3435 AVDD.n499 AVDD.n498 0.0525345
R3436 AVDD.n557 AVDD.n556 0.0525345
R3437 AVDD.n567 AVDD.n566 0.0525345
R3438 AVDD.n889 AVDD.n888 0.0525345
R3439 AVDD.n894 AVDD.n893 0.0525345
R3440 AVDD.n2142 AVDD.n2141 0.0525345
R3441 AVDD.n2148 AVDD.n2147 0.0525345
R3442 AVDD.n2161 AVDD.n2160 0.0525345
R3443 AVDD.n1059 AVDD.n1058 0.0513315
R3444 AVDD.n1006 AVDD.n744 0.0507941
R3445 AVDD.n649 AVDD.n132 0.050569
R3446 AVDD.n649 AVDD.n133 0.050569
R3447 AVDD.n1349 AVDD.n687 0.050569
R3448 AVDD.n903 AVDD.n902 0.050569
R3449 AVDD.n1349 AVDD.n1348 0.050569
R3450 AVDD.n1066 AVDD.n1065 0.0465048
R3451 AVDD.n1044 AVDD.n1043 0.0445515
R3452 AVDD.n1033 AVDD.n1032 0.0440678
R3453 AVDD.n1062 AVDD.n1061 0.0436757
R3454 AVDD.n1063 AVDD.n1062 0.0436757
R3455 AVDD.n1063 AVDD.n993 0.0436757
R3456 AVDD.n1065 AVDD.n993 0.0436757
R3457 AVDD.n1041 AVDD.n996 0.0433141
R3458 AVDD.n1040 AVDD.n996 0.0433141
R3459 AVDD.n1039 AVDD.n997 0.0433141
R3460 AVDD.n1037 AVDD.n1036 0.0433141
R3461 AVDD.n1036 AVDD.n1035 0.0433141
R3462 AVDD.n1035 AVDD.n999 0.0433141
R3463 AVDD.n1033 AVDD.n999 0.0433141
R3464 AVDD.n1042 AVDD.n1041 0.0430669
R3465 AVDD.n1179 AVDD.n1178 0.0430647
R3466 AVDD.n1131 AVDD.n751 0.0428653
R3467 AVDD.n742 AVDD.n741 0.0417941
R3468 AVDD.n1009 AVDD.n1008 0.0417941
R3469 AVDD.n604 AVDD.n603 0.0417245
R3470 AVDD.n1203 AVDD.n1202 0.0416007
R3471 AVDD.n1222 AVDD.n715 0.0415824
R3472 AVDD.n1205 AVDD.n1204 0.0413899
R3473 AVDD.n1245 AVDD.n1244 0.041314
R3474 AVDD.n1302 AVDD.n1301 0.041314
R3475 AVDD.n803 AVDD.n802 0.041314
R3476 AVDD.n1238 AVDD.n1237 0.041314
R3477 AVDD.n1297 AVDD.n1296 0.041314
R3478 AVDD.n1292 AVDD.n1291 0.041314
R3479 AVDD.n1311 AVDD.n1310 0.041314
R3480 AVDD.n806 AVDD.n805 0.041314
R3481 AVDD.n1040 AVDD.n1039 0.040902
R3482 AVDD.n366 AVDD.n365 0.0402959
R3483 AVDD.n372 AVDD.n371 0.0402959
R3484 AVDD.n399 AVDD.n398 0.0402959
R3485 AVDD.n405 AVDD.n404 0.0402959
R3486 AVDD.n612 AVDD.n611 0.0402959
R3487 AVDD.n516 AVDD.n515 0.0402959
R3488 AVDD.n519 AVDD.n518 0.0402959
R3489 AVDD.n602 AVDD.n601 0.0402959
R3490 AVDD.n1234 AVDD.n1233 0.0395167
R3491 AVDD.n1096 AVDD.n1095 0.0394276
R3492 AVDD.n598 AVDD.n597 0.0393731
R3493 AVDD.n1949 AVDD.n60 0.0392688
R3494 AVDD.n362 AVDD.n361 0.0391565
R3495 AVDD.n1011 AVDD.n1010 0.0387235
R3496 AVDD.n1098 AVDD.n982 0.0383
R3497 AVDD.n1011 AVDD.n1007 0.0373471
R3498 AVDD.n1181 AVDD.n1180 0.0371353
R3499 AVDD.n1200 AVDD.n717 0.0369637
R3500 AVDD.n1181 AVDD.n743 0.0369235
R3501 AVDD.n1201 AVDD.n1200 0.0367529
R3502 AVDD.n1494 AVDD.n1493 0.0360345
R3503 AVDD.n1498 AVDD.n111 0.0360345
R3504 AVDD.n495 AVDD.n494 0.0360345
R3505 AVDD.n563 AVDD.n562 0.0360345
R3506 AVDD.n885 AVDD.n884 0.0360345
R3507 AVDD.n899 AVDD.n898 0.0360345
R3508 AVDD.n2152 AVDD.n2151 0.0360345
R3509 AVDD.n2156 AVDD.n34 0.0360345
R3510 AVDD.n1130 AVDD.n752 0.0359624
R3511 AVDD.n2139 AVDD.n42 0.0347688
R3512 AVDD.n1538 AVDD.n87 0.0347688
R3513 AVDD.n1068 AVDD.n1067 0.0347688
R3514 AVDD.n1730 AVDD.n1729 0.0347688
R3515 AVDD.n2139 AVDD.n2138 0.0347688
R3516 AVDD.n157 AVDD.n87 0.0347688
R3517 AVDD.n1729 AVDD.n1727 0.0347688
R3518 AVDD.n369 AVDD.n368 0.0345816
R3519 AVDD.n66 AVDD.n42 0.0341759
R3520 AVDD.n1924 AVDD.n65 0.0341759
R3521 AVDD.n1927 AVDD.n65 0.0341759
R3522 AVDD.n1928 AVDD.n1927 0.0341759
R3523 AVDD.n1929 AVDD.n1928 0.0341759
R3524 AVDD.n1929 AVDD.n64 0.0341759
R3525 AVDD.n1931 AVDD.n64 0.0341759
R3526 AVDD.n1932 AVDD.n63 0.0341759
R3527 AVDD.n1934 AVDD.n63 0.0341759
R3528 AVDD.n1937 AVDD.n1936 0.0341759
R3529 AVDD.n1937 AVDD.n62 0.0341759
R3530 AVDD.n1939 AVDD.n62 0.0341759
R3531 AVDD.n1941 AVDD.n1940 0.0341759
R3532 AVDD.n1942 AVDD.n1941 0.0341759
R3533 AVDD.n1942 AVDD.n61 0.0341759
R3534 AVDD.n1945 AVDD.n61 0.0341759
R3535 AVDD.n1946 AVDD.n1945 0.0341759
R3536 AVDD.n1947 AVDD.n1946 0.0341759
R3537 AVDD.n361 AVDD.n150 0.0341759
R3538 AVDD.n359 AVDD.n358 0.0341759
R3539 AVDD.n358 AVDD.n357 0.0341759
R3540 AVDD.n357 AVDD.n348 0.0341759
R3541 AVDD.n354 AVDD.n348 0.0341759
R3542 AVDD.n354 AVDD.n353 0.0341759
R3543 AVDD.n353 AVDD.n352 0.0341759
R3544 AVDD.n351 AVDD.n349 0.0341759
R3545 AVDD.n349 AVDD.n90 0.0341759
R3546 AVDD.n1526 AVDD.n1525 0.0341759
R3547 AVDD.n1526 AVDD.n89 0.0341759
R3548 AVDD.n1528 AVDD.n89 0.0341759
R3549 AVDD.n1530 AVDD.n1529 0.0341759
R3550 AVDD.n1531 AVDD.n1530 0.0341759
R3551 AVDD.n1531 AVDD.n88 0.0341759
R3552 AVDD.n1534 AVDD.n88 0.0341759
R3553 AVDD.n1535 AVDD.n1534 0.0341759
R3554 AVDD.n1536 AVDD.n1535 0.0341759
R3555 AVDD.n1069 AVDD.n1068 0.0341759
R3556 AVDD.n1070 AVDD.n1069 0.0341759
R3557 AVDD.n1070 AVDD.n988 0.0341759
R3558 AVDD.n1073 AVDD.n988 0.0341759
R3559 AVDD.n1074 AVDD.n1073 0.0341759
R3560 AVDD.n1075 AVDD.n1074 0.0341759
R3561 AVDD.n1075 AVDD.n987 0.0341759
R3562 AVDD.n1077 AVDD.n987 0.0341759
R3563 AVDD.n1078 AVDD.n986 0.0341759
R3564 AVDD.n1080 AVDD.n986 0.0341759
R3565 AVDD.n1083 AVDD.n1082 0.0341759
R3566 AVDD.n1083 AVDD.n985 0.0341759
R3567 AVDD.n1085 AVDD.n985 0.0341759
R3568 AVDD.n1087 AVDD.n1086 0.0341759
R3569 AVDD.n1088 AVDD.n1087 0.0341759
R3570 AVDD.n1088 AVDD.n984 0.0341759
R3571 AVDD.n1091 AVDD.n984 0.0341759
R3572 AVDD.n1092 AVDD.n1091 0.0341759
R3573 AVDD.n1093 AVDD.n1092 0.0341759
R3574 AVDD.n1093 AVDD.n983 0.0341759
R3575 AVDD.n1095 AVDD.n983 0.0341759
R3576 AVDD.n1730 AVDD.n68 0.0341759
R3577 AVDD.n1756 AVDD.n69 0.0341759
R3578 AVDD.n1753 AVDD.n69 0.0341759
R3579 AVDD.n1753 AVDD.n1752 0.0341759
R3580 AVDD.n1752 AVDD.n1751 0.0341759
R3581 AVDD.n1751 AVDD.n1731 0.0341759
R3582 AVDD.n1749 AVDD.n1731 0.0341759
R3583 AVDD.n1748 AVDD.n1732 0.0341759
R3584 AVDD.n1746 AVDD.n1732 0.0341759
R3585 AVDD.n1744 AVDD.n1743 0.0341759
R3586 AVDD.n1743 AVDD.n1733 0.0341759
R3587 AVDD.n1741 AVDD.n1733 0.0341759
R3588 AVDD.n1740 AVDD.n1734 0.0341759
R3589 AVDD.n1738 AVDD.n1734 0.0341759
R3590 AVDD.n1738 AVDD.n1737 0.0341759
R3591 AVDD.n1737 AVDD.n1736 0.0341759
R3592 AVDD.n1736 AVDD.n44 0.0341759
R3593 AVDD.n2136 AVDD.n44 0.0341759
R3594 AVDD.n157 AVDD.n155 0.0341759
R3595 AVDD.n183 AVDD.n156 0.0341759
R3596 AVDD.n180 AVDD.n156 0.0341759
R3597 AVDD.n180 AVDD.n179 0.0341759
R3598 AVDD.n179 AVDD.n178 0.0341759
R3599 AVDD.n178 AVDD.n158 0.0341759
R3600 AVDD.n176 AVDD.n158 0.0341759
R3601 AVDD.n175 AVDD.n159 0.0341759
R3602 AVDD.n173 AVDD.n159 0.0341759
R3603 AVDD.n171 AVDD.n170 0.0341759
R3604 AVDD.n170 AVDD.n160 0.0341759
R3605 AVDD.n168 AVDD.n160 0.0341759
R3606 AVDD.n167 AVDD.n161 0.0341759
R3607 AVDD.n165 AVDD.n161 0.0341759
R3608 AVDD.n165 AVDD.n164 0.0341759
R3609 AVDD.n164 AVDD.n163 0.0341759
R3610 AVDD.n163 AVDD.n71 0.0341759
R3611 AVDD.n1725 AVDD.n71 0.0341759
R3612 AVDD.n569 AVDD.n448 0.0337609
R3613 AVDD.n2196 AVDD.n15 0.0337609
R3614 AVDD.n570 AVDD.n569 0.0337609
R3615 AVDD.n2196 AVDD.n2195 0.0337609
R3616 AVDD.n448 AVDD.n416 0.0331854
R3617 AVDD.n446 AVDD.n416 0.0331854
R3618 AVDD.n446 AVDD.n445 0.0331854
R3619 AVDD.n445 AVDD.n444 0.0331854
R3620 AVDD.n444 AVDD.n417 0.0331854
R3621 AVDD.n441 AVDD.n417 0.0331854
R3622 AVDD.n441 AVDD.n440 0.0331854
R3623 AVDD.n440 AVDD.n439 0.0331854
R3624 AVDD.n438 AVDD.n418 0.0331854
R3625 AVDD.n436 AVDD.n418 0.0331854
R3626 AVDD.n434 AVDD.n433 0.0331854
R3627 AVDD.n433 AVDD.n419 0.0331854
R3628 AVDD.n431 AVDD.n419 0.0331854
R3629 AVDD.n430 AVDD.n420 0.0331854
R3630 AVDD.n428 AVDD.n420 0.0331854
R3631 AVDD.n428 AVDD.n427 0.0331854
R3632 AVDD.n427 AVDD.n426 0.0331854
R3633 AVDD.n426 AVDD.n421 0.0331854
R3634 AVDD.n423 AVDD.n421 0.0331854
R3635 AVDD.n423 AVDD.n422 0.0331854
R3636 AVDD.n422 AVDD.n15 0.0331854
R3637 AVDD.n597 AVDD.n410 0.0331854
R3638 AVDD.n595 AVDD.n410 0.0331854
R3639 AVDD.n595 AVDD.n594 0.0331854
R3640 AVDD.n594 AVDD.n593 0.0331854
R3641 AVDD.n593 AVDD.n411 0.0331854
R3642 AVDD.n590 AVDD.n411 0.0331854
R3643 AVDD.n590 AVDD.n589 0.0331854
R3644 AVDD.n589 AVDD.n588 0.0331854
R3645 AVDD.n587 AVDD.n412 0.0331854
R3646 AVDD.n585 AVDD.n412 0.0331854
R3647 AVDD.n583 AVDD.n582 0.0331854
R3648 AVDD.n582 AVDD.n413 0.0331854
R3649 AVDD.n580 AVDD.n413 0.0331854
R3650 AVDD.n579 AVDD.n414 0.0331854
R3651 AVDD.n577 AVDD.n414 0.0331854
R3652 AVDD.n577 AVDD.n576 0.0331854
R3653 AVDD.n576 AVDD.n575 0.0331854
R3654 AVDD.n575 AVDD.n415 0.0331854
R3655 AVDD.n572 AVDD.n415 0.0331854
R3656 AVDD.n572 AVDD.n571 0.0331854
R3657 AVDD.n571 AVDD.n570 0.0331854
R3658 AVDD.n1231 AVDD.n1230 0.0331854
R3659 AVDD.n1231 AVDD.n712 0.0331854
R3660 AVDD.n1233 AVDD.n712 0.0331854
R3661 AVDD.n2195 AVDD.n16 0.0331854
R3662 AVDD.n2193 AVDD.n16 0.0331854
R3663 AVDD.n2193 AVDD.n2192 0.0331854
R3664 AVDD.n2192 AVDD.n2191 0.0331854
R3665 AVDD.n2191 AVDD.n17 0.0331854
R3666 AVDD.n2188 AVDD.n17 0.0331854
R3667 AVDD.n2188 AVDD.n2187 0.0331854
R3668 AVDD.n2187 AVDD.n2186 0.0331854
R3669 AVDD.n2185 AVDD.n18 0.0331854
R3670 AVDD.n2183 AVDD.n18 0.0331854
R3671 AVDD.n909 AVDD.n19 0.0331854
R3672 AVDD.n909 AVDD.n908 0.0331854
R3673 AVDD.n911 AVDD.n908 0.0331854
R3674 AVDD.n912 AVDD.n907 0.0331854
R3675 AVDD.n914 AVDD.n907 0.0331854
R3676 AVDD.n915 AVDD.n914 0.0331854
R3677 AVDD.n918 AVDD.n915 0.0331854
R3678 AVDD.n1932 AVDD.n1931 0.0325158
R3679 AVDD.n1940 AVDD.n1939 0.0325158
R3680 AVDD.n352 AVDD.n351 0.0325158
R3681 AVDD.n1529 AVDD.n1528 0.0325158
R3682 AVDD.n1078 AVDD.n1077 0.0325158
R3683 AVDD.n1086 AVDD.n1085 0.0325158
R3684 AVDD.n1749 AVDD.n1748 0.0325158
R3685 AVDD.n1741 AVDD.n1740 0.0325158
R3686 AVDD.n176 AVDD.n175 0.0325158
R3687 AVDD.n168 AVDD.n167 0.0325158
R3688 AVDD.n741 AVDD.n715 0.0320529
R3689 AVDD.n743 AVDD.n742 0.0320529
R3690 AVDD.n1180 AVDD.n1179 0.0320529
R3691 AVDD.n1007 AVDD.n1006 0.0320529
R3692 AVDD.n1010 AVDD.n1009 0.0320529
R3693 AVDD.n1008 AVDD.n982 0.0320529
R3694 AVDD.n1097 AVDD.n1096 0.0320529
R3695 AVDD.n1464 AVDD.n1458 0.0319413
R3696 AVDD.n1464 AVDD.n1463 0.0319104
R3697 AVDD.n1204 AVDD.n1203 0.0319052
R3698 AVDD.n1202 AVDD.n1201 0.0319052
R3699 AVDD.n751 AVDD.n717 0.0319052
R3700 AVDD.n1242 AVDD.n60 0.031686
R3701 AVDD.n1244 AVDD.n1243 0.031686
R3702 AVDD.n1246 AVDD.n1245 0.031686
R3703 AVDD.n1303 AVDD.n1302 0.031686
R3704 AVDD.n1301 AVDD.n1300 0.031686
R3705 AVDD.n804 AVDD.n803 0.031686
R3706 AVDD.n802 AVDD.n711 0.031686
R3707 AVDD.n1239 AVDD.n1238 0.031686
R3708 AVDD.n1237 AVDD.n1236 0.031686
R3709 AVDD.n1235 AVDD.n1234 0.031686
R3710 AVDD.n1298 AVDD.n1297 0.031686
R3711 AVDD.n1296 AVDD.n1295 0.031686
R3712 AVDD.n1293 AVDD.n1292 0.031686
R3713 AVDD.n1291 AVDD.n705 0.031686
R3714 AVDD.n1312 AVDD.n1311 0.031686
R3715 AVDD.n1310 AVDD.n1309 0.031686
R3716 AVDD.n805 AVDD.n706 0.031686
R3717 AVDD.n807 AVDD.n806 0.031686
R3718 AVDD.n439 AVDD.n438 0.0315742
R3719 AVDD.n431 AVDD.n430 0.0315742
R3720 AVDD.n588 AVDD.n587 0.0315742
R3721 AVDD.n580 AVDD.n579 0.0315742
R3722 AVDD.n2186 AVDD.n2185 0.0315742
R3723 AVDD.n912 AVDD.n911 0.0315742
R3724 AVDD.n1442 AVDD.n1441 0.0315707
R3725 AVDD.n1447 AVDD.n1446 0.0315707
R3726 AVDD.n1457 AVDD.n1456 0.0315707
R3727 AVDD.n1462 AVDD.n1461 0.0315707
R3728 AVDD.n2213 AVDD.n2212 0.0315707
R3729 AVDD.n2208 AVDD.n2207 0.0315707
R3730 AVDD.n2199 AVDD.n2198 0.0315707
R3731 AVDD.n1494 AVDD.n1488 0.0313793
R3732 AVDD.n1499 AVDD.n1498 0.0313793
R3733 AVDD.n494 AVDD.n492 0.0313793
R3734 AVDD.n562 AVDD.n560 0.0313793
R3735 AVDD.n884 AVDD.n882 0.0313793
R3736 AVDD.n898 AVDD.n897 0.0313793
R3737 AVDD.n2152 AVDD.n2145 0.0313793
R3738 AVDD.n2157 AVDD.n2156 0.0313793
R3739 AVDD.n1230 AVDD.n1229 0.0311937
R3740 AVDD.n363 AVDD.n362 0.0309082
R3741 AVDD.n365 AVDD.n364 0.0309082
R3742 AVDD.n367 AVDD.n366 0.0309082
R3743 AVDD.n371 AVDD.n370 0.0309082
R3744 AVDD.n373 AVDD.n372 0.0309082
R3745 AVDD.n398 AVDD.n397 0.0309082
R3746 AVDD.n400 AVDD.n399 0.0309082
R3747 AVDD.n404 AVDD.n403 0.0309082
R3748 AVDD.n406 AVDD.n405 0.0309082
R3749 AVDD.n613 AVDD.n612 0.0309082
R3750 AVDD.n611 AVDD.n610 0.0309082
R3751 AVDD.n515 AVDD.n514 0.0309082
R3752 AVDD.n517 AVDD.n516 0.0309082
R3753 AVDD.n520 AVDD.n519 0.0309082
R3754 AVDD.n518 AVDD.n408 0.0309082
R3755 AVDD.n603 AVDD.n602 0.0309082
R3756 AVDD.n601 AVDD.n600 0.0309082
R3757 AVDD.n599 AVDD.n598 0.0309082
R3758 AVDD.n1935 AVDD.n1934 0.0303814
R3759 AVDD.n1524 AVDD.n90 0.0303814
R3760 AVDD.n1746 AVDD.n1745 0.0303814
R3761 AVDD.n173 AVDD.n172 0.0303814
R3762 AVDD.n1950 AVDD.n1949 0.0302628
R3763 AVDD.n1539 AVDD.n1538 0.0302628
R3764 AVDD.n2138 AVDD.n43 0.0302628
R3765 AVDD.n1727 AVDD.n70 0.0302628
R3766 AVDD.n1081 AVDD.n1080 0.0295514
R3767 AVDD.n436 AVDD.n435 0.0295026
R3768 AVDD.n585 AVDD.n584 0.0295026
R3769 AVDD.n2183 AVDD.n2182 0.0295026
R3770 AVDD.n605 AVDD.n604 0.0293776
R3771 AVDD.n1046 AVDD.n1045 0.0289485
R3772 AVDD.n368 AVDD.n367 0.0273367
R3773 AVDD.n1058 AVDD.n994 0.0261926
R3774 AVDD.n998 AVDD.n997 0.0259774
R3775 AVDD.n1043 AVDD.n1042 0.0234742
R3776 AVDD.n1045 AVDD.n1044 0.0234742
R3777 AVDD.n1505 AVDD.n110 0.0228966
R3778 AVDD.n554 AVDD.n500 0.0228966
R3779 AVDD.n891 AVDD.n890 0.0228966
R3780 AVDD.n2163 AVDD.n33 0.0228966
R3781 AVDD.n1505 AVDD.n1504 0.0228448
R3782 AVDD.n555 AVDD.n554 0.0228448
R3783 AVDD.n892 AVDD.n891 0.0228448
R3784 AVDD.n2163 AVDD.n2162 0.0228448
R3785 AVDD.n1055 AVDD.n1054 0.0224615
R3786 AVDD.n2221 AVDD.n2 0.0217183
R3787 AVDD.n1453 AVDD.n1452 0.0217183
R3788 AVDD.n2217 AVDD.n2216 0.0217183
R3789 AVDD.n2203 AVDD.n2202 0.0217183
R3790 AVDD.n1487 AVDD.n1486 0.0206724
R3791 AVDD.n1492 AVDD.n1491 0.0206724
R3792 AVDD.n1501 AVDD.n1500 0.0206724
R3793 AVDD.n131 AVDD.n130 0.0206724
R3794 AVDD.n491 AVDD.n490 0.0206724
R3795 AVDD.n497 AVDD.n496 0.0206724
R3796 AVDD.n559 AVDD.n558 0.0206724
R3797 AVDD.n565 AVDD.n564 0.0206724
R3798 AVDD.n881 AVDD.n880 0.0206724
R3799 AVDD.n887 AVDD.n886 0.0206724
R3800 AVDD.n896 AVDD.n895 0.0206724
R3801 AVDD.n901 AVDD.n900 0.0206724
R3802 AVDD.n2144 AVDD.n2143 0.0206724
R3803 AVDD.n2150 AVDD.n2149 0.0206724
R3804 AVDD.n2159 AVDD.n2158 0.0206724
R3805 AVDD.n1347 AVDD.n1346 0.0206724
R3806 AVDD.n1947 AVDD.n58 0.0204161
R3807 AVDD.n1536 AVDD.n85 0.0204161
R3808 AVDD.n2136 AVDD.n2135 0.0204161
R3809 AVDD.n1725 AVDD.n1724 0.0204161
R3810 AVDD.n1923 AVDD.n66 0.019782
R3811 AVDD.n347 AVDD.n150 0.019782
R3812 AVDD.n1757 AVDD.n68 0.019782
R3813 AVDD.n184 AVDD.n155 0.019782
R3814 AVDD.n394 AVDD.n393 0.0196477
R3815 AVDD.n524 AVDD.n523 0.0196477
R3816 AVDD.n811 AVDD.n810 0.0196477
R3817 AVDD.n1289 AVDD.n1288 0.0196477
R3818 AVDD.n2222 AVDD.n2221 0.0189386
R3819 AVDD.n1452 AVDD.n1450 0.0189386
R3820 AVDD.n2217 AVDD.n10 0.0189386
R3821 AVDD.n2204 AVDD.n2203 0.0189386
R3822 AVDD.n1029 AVDD.n1028 0.0185
R3823 AVDD AVDD.n2225 0.0182591
R3824 AVDD.n1061 AVDD.n994 0.0179831
R3825 AVDD.n1037 AVDD.n998 0.0178367
R3826 AVDD.n1924 AVDD.n1923 0.0177463
R3827 AVDD.n359 AVDD.n347 0.0177463
R3828 AVDD.n1757 AVDD.n1756 0.0177463
R3829 AVDD.n184 AVDD.n183 0.0177463
R3830 AVDD.n1444 AVDD.n1398 0.0174226
R3831 AVDD.n2164 AVDD.n2163 0.0174226
R3832 AVDD.n554 AVDD.n489 0.0174226
R3833 AVDD.n2210 AVDD.n12 0.0174226
R3834 AVDD.n1505 AVDD.n109 0.0174226
R3835 AVDD.n1444 AVDD.n1438 0.0174226
R3836 AVDD.n1506 AVDD.n1505 0.0174226
R3837 AVDD.n554 AVDD.n553 0.0174226
R3838 AVDD.n891 AVDD.n838 0.0174226
R3839 AVDD.n2210 AVDD.n13 0.0174226
R3840 AVDD.n891 AVDD.n879 0.0174226
R3841 AVDD.n2163 AVDD.n32 0.0174226
R3842 AVDD.n1398 AVDD.n1380 0.0171298
R3843 AVDD.n1396 AVDD.n1380 0.0171298
R3844 AVDD.n1396 AVDD.n1395 0.0171298
R3845 AVDD.n1395 AVDD.n1394 0.0171298
R3846 AVDD.n1394 AVDD.n1383 0.0171298
R3847 AVDD.n1391 AVDD.n1383 0.0171298
R3848 AVDD.n1391 AVDD.n1390 0.0171298
R3849 AVDD.n1390 AVDD.n1389 0.0171298
R3850 AVDD.n1388 AVDD.n1386 0.0171298
R3851 AVDD.n1386 AVDD.n24 0.0171298
R3852 AVDD.n2177 AVDD.n2176 0.0171298
R3853 AVDD.n2176 AVDD.n26 0.0171298
R3854 AVDD.n2174 AVDD.n26 0.0171298
R3855 AVDD.n2173 AVDD.n27 0.0171298
R3856 AVDD.n2171 AVDD.n27 0.0171298
R3857 AVDD.n2171 AVDD.n2170 0.0171298
R3858 AVDD.n2170 AVDD.n2169 0.0171298
R3859 AVDD.n2169 AVDD.n30 0.0171298
R3860 AVDD.n2166 AVDD.n30 0.0171298
R3861 AVDD.n2166 AVDD.n2165 0.0171298
R3862 AVDD.n2165 AVDD.n2164 0.0171298
R3863 AVDD.n489 AVDD.n449 0.0171298
R3864 AVDD.n487 AVDD.n449 0.0171298
R3865 AVDD.n487 AVDD.n486 0.0171298
R3866 AVDD.n486 AVDD.n485 0.0171298
R3867 AVDD.n485 AVDD.n452 0.0171298
R3868 AVDD.n482 AVDD.n452 0.0171298
R3869 AVDD.n482 AVDD.n481 0.0171298
R3870 AVDD.n481 AVDD.n480 0.0171298
R3871 AVDD.n479 AVDD.n454 0.0171298
R3872 AVDD.n477 AVDD.n454 0.0171298
R3873 AVDD.n475 AVDD.n474 0.0171298
R3874 AVDD.n474 AVDD.n457 0.0171298
R3875 AVDD.n472 AVDD.n457 0.0171298
R3876 AVDD.n471 AVDD.n458 0.0171298
R3877 AVDD.n469 AVDD.n458 0.0171298
R3878 AVDD.n469 AVDD.n468 0.0171298
R3879 AVDD.n468 AVDD.n467 0.0171298
R3880 AVDD.n467 AVDD.n461 0.0171298
R3881 AVDD.n464 AVDD.n461 0.0171298
R3882 AVDD.n464 AVDD.n463 0.0171298
R3883 AVDD.n463 AVDD.n12 0.0171298
R3884 AVDD.n1409 AVDD.n109 0.0171298
R3885 AVDD.n1411 AVDD.n1409 0.0171298
R3886 AVDD.n1411 AVDD.n1408 0.0171298
R3887 AVDD.n1414 AVDD.n1408 0.0171298
R3888 AVDD.n1414 AVDD.n1407 0.0171298
R3889 AVDD.n1417 AVDD.n1407 0.0171298
R3890 AVDD.n1417 AVDD.n1406 0.0171298
R3891 AVDD.n1419 AVDD.n1406 0.0171298
R3892 AVDD.n1420 AVDD.n1405 0.0171298
R3893 AVDD.n1422 AVDD.n1405 0.0171298
R3894 AVDD.n1425 AVDD.n1404 0.0171298
R3895 AVDD.n1425 AVDD.n1403 0.0171298
R3896 AVDD.n1427 AVDD.n1403 0.0171298
R3897 AVDD.n1428 AVDD.n1402 0.0171298
R3898 AVDD.n1430 AVDD.n1402 0.0171298
R3899 AVDD.n1430 AVDD.n1401 0.0171298
R3900 AVDD.n1433 AVDD.n1401 0.0171298
R3901 AVDD.n1433 AVDD.n1400 0.0171298
R3902 AVDD.n1436 AVDD.n1400 0.0171298
R3903 AVDD.n1436 AVDD.n1399 0.0171298
R3904 AVDD.n1438 AVDD.n1399 0.0171298
R3905 AVDD.n395 AVDD.n394 0.0171298
R3906 AVDD.n393 AVDD.n375 0.0171298
R3907 AVDD.n391 AVDD.n375 0.0171298
R3908 AVDD.n391 AVDD.n390 0.0171298
R3909 AVDD.n390 AVDD.n389 0.0171298
R3910 AVDD.n389 AVDD.n378 0.0171298
R3911 AVDD.n386 AVDD.n378 0.0171298
R3912 AVDD.n386 AVDD.n385 0.0171298
R3913 AVDD.n385 AVDD.n384 0.0171298
R3914 AVDD.n383 AVDD.n381 0.0171298
R3915 AVDD.n381 AVDD.n101 0.0171298
R3916 AVDD.n1519 AVDD.n1518 0.0171298
R3917 AVDD.n1518 AVDD.n103 0.0171298
R3918 AVDD.n1516 AVDD.n103 0.0171298
R3919 AVDD.n1515 AVDD.n104 0.0171298
R3920 AVDD.n1513 AVDD.n104 0.0171298
R3921 AVDD.n1513 AVDD.n1512 0.0171298
R3922 AVDD.n1512 AVDD.n1511 0.0171298
R3923 AVDD.n1511 AVDD.n107 0.0171298
R3924 AVDD.n1508 AVDD.n107 0.0171298
R3925 AVDD.n1508 AVDD.n1507 0.0171298
R3926 AVDD.n1507 AVDD.n1506 0.0171298
R3927 AVDD.n523 AVDD.n513 0.0171298
R3928 AVDD.n524 AVDD.n512 0.0171298
R3929 AVDD.n526 AVDD.n512 0.0171298
R3930 AVDD.n526 AVDD.n511 0.0171298
R3931 AVDD.n529 AVDD.n511 0.0171298
R3932 AVDD.n529 AVDD.n510 0.0171298
R3933 AVDD.n532 AVDD.n510 0.0171298
R3934 AVDD.n532 AVDD.n509 0.0171298
R3935 AVDD.n534 AVDD.n509 0.0171298
R3936 AVDD.n535 AVDD.n507 0.0171298
R3937 AVDD.n537 AVDD.n507 0.0171298
R3938 AVDD.n540 AVDD.n506 0.0171298
R3939 AVDD.n540 AVDD.n505 0.0171298
R3940 AVDD.n542 AVDD.n505 0.0171298
R3941 AVDD.n543 AVDD.n504 0.0171298
R3942 AVDD.n545 AVDD.n504 0.0171298
R3943 AVDD.n545 AVDD.n503 0.0171298
R3944 AVDD.n548 AVDD.n503 0.0171298
R3945 AVDD.n548 AVDD.n502 0.0171298
R3946 AVDD.n551 AVDD.n502 0.0171298
R3947 AVDD.n551 AVDD.n501 0.0171298
R3948 AVDD.n553 AVDD.n501 0.0171298
R3949 AVDD.n838 AVDD.n787 0.0171298
R3950 AVDD.n836 AVDD.n787 0.0171298
R3951 AVDD.n836 AVDD.n835 0.0171298
R3952 AVDD.n835 AVDD.n834 0.0171298
R3953 AVDD.n834 AVDD.n790 0.0171298
R3954 AVDD.n831 AVDD.n790 0.0171298
R3955 AVDD.n831 AVDD.n830 0.0171298
R3956 AVDD.n830 AVDD.n829 0.0171298
R3957 AVDD.n828 AVDD.n792 0.0171298
R3958 AVDD.n826 AVDD.n792 0.0171298
R3959 AVDD.n824 AVDD.n823 0.0171298
R3960 AVDD.n823 AVDD.n795 0.0171298
R3961 AVDD.n821 AVDD.n795 0.0171298
R3962 AVDD.n820 AVDD.n796 0.0171298
R3963 AVDD.n818 AVDD.n796 0.0171298
R3964 AVDD.n818 AVDD.n817 0.0171298
R3965 AVDD.n817 AVDD.n816 0.0171298
R3966 AVDD.n816 AVDD.n799 0.0171298
R3967 AVDD.n813 AVDD.n799 0.0171298
R3968 AVDD.n813 AVDD.n812 0.0171298
R3969 AVDD.n812 AVDD.n811 0.0171298
R3970 AVDD.n810 AVDD.n801 0.0171298
R3971 AVDD.n850 AVDD.n13 0.0171298
R3972 AVDD.n852 AVDD.n850 0.0171298
R3973 AVDD.n852 AVDD.n849 0.0171298
R3974 AVDD.n855 AVDD.n849 0.0171298
R3975 AVDD.n855 AVDD.n848 0.0171298
R3976 AVDD.n858 AVDD.n848 0.0171298
R3977 AVDD.n858 AVDD.n847 0.0171298
R3978 AVDD.n860 AVDD.n847 0.0171298
R3979 AVDD.n861 AVDD.n845 0.0171298
R3980 AVDD.n863 AVDD.n845 0.0171298
R3981 AVDD.n866 AVDD.n844 0.0171298
R3982 AVDD.n866 AVDD.n843 0.0171298
R3983 AVDD.n868 AVDD.n843 0.0171298
R3984 AVDD.n869 AVDD.n842 0.0171298
R3985 AVDD.n871 AVDD.n842 0.0171298
R3986 AVDD.n871 AVDD.n841 0.0171298
R3987 AVDD.n874 AVDD.n841 0.0171298
R3988 AVDD.n874 AVDD.n840 0.0171298
R3989 AVDD.n877 AVDD.n840 0.0171298
R3990 AVDD.n877 AVDD.n839 0.0171298
R3991 AVDD.n879 AVDD.n839 0.0171298
R3992 AVDD.n1259 AVDD.n32 0.0171298
R3993 AVDD.n1261 AVDD.n1259 0.0171298
R3994 AVDD.n1261 AVDD.n1258 0.0171298
R3995 AVDD.n1264 AVDD.n1258 0.0171298
R3996 AVDD.n1264 AVDD.n1257 0.0171298
R3997 AVDD.n1267 AVDD.n1257 0.0171298
R3998 AVDD.n1267 AVDD.n1256 0.0171298
R3999 AVDD.n1269 AVDD.n1256 0.0171298
R4000 AVDD.n1270 AVDD.n1254 0.0171298
R4001 AVDD.n1272 AVDD.n1254 0.0171298
R4002 AVDD.n1275 AVDD.n1253 0.0171298
R4003 AVDD.n1275 AVDD.n1252 0.0171298
R4004 AVDD.n1277 AVDD.n1252 0.0171298
R4005 AVDD.n1278 AVDD.n1251 0.0171298
R4006 AVDD.n1280 AVDD.n1251 0.0171298
R4007 AVDD.n1280 AVDD.n1250 0.0171298
R4008 AVDD.n1283 AVDD.n1250 0.0171298
R4009 AVDD.n1283 AVDD.n1249 0.0171298
R4010 AVDD.n1286 AVDD.n1249 0.0171298
R4011 AVDD.n1286 AVDD.n1248 0.0171298
R4012 AVDD.n1288 AVDD.n1248 0.0171298
R4013 AVDD.n1289 AVDD.n1247 0.0171298
R4014 AVDD.n374 AVDD.n149 0.0166614
R4015 AVDD.n522 AVDD.n409 0.0166614
R4016 AVDD.n1051 AVDD.n1050 0.0163144
R4017 AVDD.n1389 AVDD.n1388 0.01631
R4018 AVDD.n2174 AVDD.n2173 0.01631
R4019 AVDD.n480 AVDD.n479 0.01631
R4020 AVDD.n472 AVDD.n471 0.01631
R4021 AVDD.n1420 AVDD.n1419 0.01631
R4022 AVDD.n1428 AVDD.n1427 0.01631
R4023 AVDD.n384 AVDD.n383 0.01631
R4024 AVDD.n1516 AVDD.n1515 0.01631
R4025 AVDD.n535 AVDD.n534 0.01631
R4026 AVDD.n543 AVDD.n542 0.01631
R4027 AVDD.n829 AVDD.n828 0.01631
R4028 AVDD.n821 AVDD.n820 0.01631
R4029 AVDD.n861 AVDD.n860 0.01631
R4030 AVDD.n869 AVDD.n868 0.01631
R4031 AVDD.n1270 AVDD.n1269 0.01631
R4032 AVDD.n1278 AVDD.n1277 0.01631
R4033 AVDD.n59 AVDD.n58 0.0162238
R4034 AVDD.n86 AVDD.n85 0.0162238
R4035 AVDD.n2135 AVDD.n45 0.0162238
R4036 AVDD.n1724 AVDD.n72 0.0162238
R4037 AVDD.n1484 AVDD.n1483 0.0159138
R4038 AVDD.n1486 AVDD.n1485 0.0159138
R4039 AVDD.n1488 AVDD.n1487 0.0159138
R4040 AVDD.n1493 AVDD.n1492 0.0159138
R4041 AVDD.n1491 AVDD.n1490 0.0159138
R4042 AVDD.n1489 AVDD.n110 0.0159138
R4043 AVDD.n1504 AVDD.n1503 0.0159138
R4044 AVDD.n1502 AVDD.n1501 0.0159138
R4045 AVDD.n1500 AVDD.n1499 0.0159138
R4046 AVDD.n130 AVDD.n111 0.0159138
R4047 AVDD.n132 AVDD.n131 0.0159138
R4048 AVDD.n490 AVDD.n133 0.0159138
R4049 AVDD.n492 AVDD.n491 0.0159138
R4050 AVDD.n496 AVDD.n495 0.0159138
R4051 AVDD.n498 AVDD.n497 0.0159138
R4052 AVDD.n500 AVDD.n499 0.0159138
R4053 AVDD.n556 AVDD.n555 0.0159138
R4054 AVDD.n558 AVDD.n557 0.0159138
R4055 AVDD.n560 AVDD.n559 0.0159138
R4056 AVDD.n564 AVDD.n563 0.0159138
R4057 AVDD.n566 AVDD.n565 0.0159138
R4058 AVDD.n568 AVDD.n567 0.0159138
R4059 AVDD.n880 AVDD.n687 0.0159138
R4060 AVDD.n882 AVDD.n881 0.0159138
R4061 AVDD.n886 AVDD.n885 0.0159138
R4062 AVDD.n888 AVDD.n887 0.0159138
R4063 AVDD.n890 AVDD.n889 0.0159138
R4064 AVDD.n893 AVDD.n892 0.0159138
R4065 AVDD.n895 AVDD.n894 0.0159138
R4066 AVDD.n897 AVDD.n896 0.0159138
R4067 AVDD.n900 AVDD.n899 0.0159138
R4068 AVDD.n902 AVDD.n901 0.0159138
R4069 AVDD.n2141 AVDD.n2140 0.0159138
R4070 AVDD.n2143 AVDD.n2142 0.0159138
R4071 AVDD.n2145 AVDD.n2144 0.0159138
R4072 AVDD.n2151 AVDD.n2150 0.0159138
R4073 AVDD.n2149 AVDD.n2148 0.0159138
R4074 AVDD.n2147 AVDD.n33 0.0159138
R4075 AVDD.n2162 AVDD.n2161 0.0159138
R4076 AVDD.n2160 AVDD.n2159 0.0159138
R4077 AVDD.n2158 AVDD.n2157 0.0159138
R4078 AVDD.n1346 AVDD.n34 0.0159138
R4079 AVDD.n1348 AVDD.n1347 0.0159138
R4080 AVDD.n1053 AVDD.n1052 0.0156839
R4081 AVDD.n1050 AVDD.n1047 0.0154737
R4082 AVDD.n2178 AVDD.n24 0.015256
R4083 AVDD.n477 AVDD.n476 0.015256
R4084 AVDD.n1422 AVDD.n118 0.015256
R4085 AVDD.n1520 AVDD.n101 0.015256
R4086 AVDD.n537 AVDD.n508 0.015256
R4087 AVDD.n826 AVDD.n825 0.015256
R4088 AVDD.n863 AVDD.n846 0.015256
R4089 AVDD.n1272 AVDD.n1255 0.015256
R4090 AVDD.n1121 AVDD.n1120 0.0148793
R4091 AVDD.n1000 AVDD.n957 0.0142069
R4092 AVDD.n1444 AVDD.n1443 0.0138734
R4093 AVDD.n2211 AVDD.n2210 0.0138734
R4094 AVDD.n990 AVDD.n989 0.0138448
R4095 AVDD.n1445 AVDD.n1444 0.0138425
R4096 AVDD.n2210 AVDD.n2209 0.0138425
R4097 AVDD AVDD.n0 0.0138116
R4098 AVDD.n918 AVDD.n917 0.012725
R4099 AVDD.n2224 AVDD.n2223 0.0125453
R4100 AVDD.n1440 AVDD.n1439 0.0125453
R4101 AVDD.n1449 AVDD.n1448 0.0125453
R4102 AVDD.n1455 AVDD.n1454 0.0125453
R4103 AVDD.n1460 AVDD.n1459 0.0125453
R4104 AVDD.n2215 AVDD.n2214 0.0125453
R4105 AVDD.n2206 AVDD.n2205 0.0125453
R4106 AVDD.n2201 AVDD.n2200 0.0125453
R4107 AVDD.n1047 AVDD.n1046 0.0119536
R4108 AVDD.n1052 AVDD.n1051 0.0119536
R4109 AVDD.n1054 AVDD.n1053 0.0119536
R4110 AVDD.n1031 AVDD.n1030 0.0117759
R4111 AVDD.n1005 AVDD.n1004 0.0117759
R4112 AVDD.n1119 AVDD.n1118 0.0117759
R4113 AVDD.n989 AVDD.n958 0.0117759
R4114 AVDD.n1057 AVDD.n1056 0.0116909
R4115 AVDD.n617 AVDD.n616 0.0113718
R4116 AVDD.n647 AVDD.n646 0.0113718
R4117 AVDD.n652 AVDD.n651 0.0113718
R4118 AVDD.n1352 AVDD.n1351 0.0113718
R4119 AVDD.n1344 AVDD.n1343 0.0113718
R4120 AVDD.n1316 AVDD.n1315 0.0113718
R4121 AVDD.n1003 AVDD.n1002 0.0111034
R4122 AVDD.n809 AVDD.n808 0.0108058
R4123 AVDD.n1299 AVDD.n1290 0.0108058
R4124 AVDD.n396 AVDD.n374 0.0101617
R4125 AVDD.n522 AVDD.n521 0.0101617
R4126 AVDD.n1465 AVDD.n1464 0.0101084
R4127 AVDD.n1464 AVDD.n1379 0.0101084
R4128 AVDD.n616 AVDD.n147 0.00994219
R4129 AVDD.n617 AVDD.n146 0.00994219
R4130 AVDD.n619 AVDD.n146 0.00994219
R4131 AVDD.n619 AVDD.n145 0.00994219
R4132 AVDD.n622 AVDD.n145 0.00994219
R4133 AVDD.n622 AVDD.n144 0.00994219
R4134 AVDD.n625 AVDD.n144 0.00994219
R4135 AVDD.n625 AVDD.n143 0.00994219
R4136 AVDD.n627 AVDD.n143 0.00994219
R4137 AVDD.n628 AVDD.n141 0.00994219
R4138 AVDD.n630 AVDD.n141 0.00994219
R4139 AVDD.n633 AVDD.n140 0.00994219
R4140 AVDD.n633 AVDD.n139 0.00994219
R4141 AVDD.n635 AVDD.n139 0.00994219
R4142 AVDD.n636 AVDD.n138 0.00994219
R4143 AVDD.n638 AVDD.n138 0.00994219
R4144 AVDD.n638 AVDD.n137 0.00994219
R4145 AVDD.n641 AVDD.n137 0.00994219
R4146 AVDD.n641 AVDD.n136 0.00994219
R4147 AVDD.n644 AVDD.n136 0.00994219
R4148 AVDD.n644 AVDD.n135 0.00994219
R4149 AVDD.n646 AVDD.n135 0.00994219
R4150 AVDD.n647 AVDD.n134 0.00994219
R4151 AVDD.n648 AVDD.n134 0.00994219
R4152 AVDD.n650 AVDD.n129 0.00994219
R4153 AVDD.n651 AVDD.n129 0.00994219
R4154 AVDD.n652 AVDD.n128 0.00994219
R4155 AVDD.n654 AVDD.n128 0.00994219
R4156 AVDD.n654 AVDD.n127 0.00994219
R4157 AVDD.n657 AVDD.n127 0.00994219
R4158 AVDD.n657 AVDD.n126 0.00994219
R4159 AVDD.n660 AVDD.n126 0.00994219
R4160 AVDD.n660 AVDD.n125 0.00994219
R4161 AVDD.n662 AVDD.n125 0.00994219
R4162 AVDD.n665 AVDD.n664 0.00994219
R4163 AVDD.n664 AVDD.n122 0.00994219
R4164 AVDD.n1478 AVDD.n1477 0.00994219
R4165 AVDD.n1477 AVDD.n124 0.00994219
R4166 AVDD.n1475 AVDD.n124 0.00994219
R4167 AVDD.n1474 AVDD.n667 0.00994219
R4168 AVDD.n1472 AVDD.n667 0.00994219
R4169 AVDD.n1472 AVDD.n1471 0.00994219
R4170 AVDD.n1471 AVDD.n1470 0.00994219
R4171 AVDD.n1470 AVDD.n670 0.00994219
R4172 AVDD.n1467 AVDD.n670 0.00994219
R4173 AVDD.n1467 AVDD.n1466 0.00994219
R4174 AVDD.n1466 AVDD.n1465 0.00994219
R4175 AVDD.n1379 AVDD.n672 0.00994219
R4176 AVDD.n1377 AVDD.n672 0.00994219
R4177 AVDD.n1377 AVDD.n1376 0.00994219
R4178 AVDD.n1376 AVDD.n1375 0.00994219
R4179 AVDD.n1375 AVDD.n675 0.00994219
R4180 AVDD.n1372 AVDD.n675 0.00994219
R4181 AVDD.n1372 AVDD.n1371 0.00994219
R4182 AVDD.n1371 AVDD.n1370 0.00994219
R4183 AVDD.n1369 AVDD.n677 0.00994219
R4184 AVDD.n1367 AVDD.n677 0.00994219
R4185 AVDD.n1365 AVDD.n1364 0.00994219
R4186 AVDD.n1364 AVDD.n680 0.00994219
R4187 AVDD.n1362 AVDD.n680 0.00994219
R4188 AVDD.n1361 AVDD.n681 0.00994219
R4189 AVDD.n1359 AVDD.n681 0.00994219
R4190 AVDD.n1359 AVDD.n1358 0.00994219
R4191 AVDD.n1358 AVDD.n1357 0.00994219
R4192 AVDD.n1357 AVDD.n684 0.00994219
R4193 AVDD.n1354 AVDD.n684 0.00994219
R4194 AVDD.n1354 AVDD.n1353 0.00994219
R4195 AVDD.n1353 AVDD.n1352 0.00994219
R4196 AVDD.n1351 AVDD.n686 0.00994219
R4197 AVDD.n1350 AVDD.n686 0.00994219
R4198 AVDD.n1345 AVDD.n688 0.00994219
R4199 AVDD.n1344 AVDD.n688 0.00994219
R4200 AVDD.n1343 AVDD.n689 0.00994219
R4201 AVDD.n1341 AVDD.n689 0.00994219
R4202 AVDD.n1341 AVDD.n1340 0.00994219
R4203 AVDD.n1340 AVDD.n1339 0.00994219
R4204 AVDD.n1339 AVDD.n692 0.00994219
R4205 AVDD.n1336 AVDD.n692 0.00994219
R4206 AVDD.n1336 AVDD.n1335 0.00994219
R4207 AVDD.n1335 AVDD.n1334 0.00994219
R4208 AVDD.n1333 AVDD.n694 0.00994219
R4209 AVDD.n1331 AVDD.n694 0.00994219
R4210 AVDD.n1329 AVDD.n1328 0.00994219
R4211 AVDD.n1328 AVDD.n698 0.00994219
R4212 AVDD.n1326 AVDD.n698 0.00994219
R4213 AVDD.n1325 AVDD.n699 0.00994219
R4214 AVDD.n1323 AVDD.n699 0.00994219
R4215 AVDD.n1323 AVDD.n1322 0.00994219
R4216 AVDD.n1322 AVDD.n1321 0.00994219
R4217 AVDD.n1321 AVDD.n702 0.00994219
R4218 AVDD.n1318 AVDD.n702 0.00994219
R4219 AVDD.n1318 AVDD.n1317 0.00994219
R4220 AVDD.n1317 AVDD.n1316 0.00994219
R4221 AVDD.n1315 AVDD.n704 0.00994219
R4222 AVDD.n1728 AVDD.n0 0.00970384
R4223 AVDD.n2225 AVDD.n2224 0.00970384
R4224 AVDD.n2223 AVDD.n2222 0.00970384
R4225 AVDD.n1439 AVDD.n2 0.00970384
R4226 AVDD.n1441 AVDD.n1440 0.00970384
R4227 AVDD.n1443 AVDD.n1442 0.00970384
R4228 AVDD.n1446 AVDD.n1445 0.00970384
R4229 AVDD.n1448 AVDD.n1447 0.00970384
R4230 AVDD.n1450 AVDD.n1449 0.00970384
R4231 AVDD.n1454 AVDD.n1453 0.00970384
R4232 AVDD.n1456 AVDD.n1455 0.00970384
R4233 AVDD.n1458 AVDD.n1457 0.00970384
R4234 AVDD.n1463 AVDD.n1462 0.00970384
R4235 AVDD.n1461 AVDD.n1460 0.00970384
R4236 AVDD.n1459 AVDD.n10 0.00970384
R4237 AVDD.n2216 AVDD.n2215 0.00970384
R4238 AVDD.n2214 AVDD.n2213 0.00970384
R4239 AVDD.n2212 AVDD.n2211 0.00970384
R4240 AVDD.n2209 AVDD.n2208 0.00970384
R4241 AVDD.n2207 AVDD.n2206 0.00970384
R4242 AVDD.n2205 AVDD.n2204 0.00970384
R4243 AVDD.n2202 AVDD.n2201 0.00970384
R4244 AVDD.n2200 AVDD.n2199 0.00970384
R4245 AVDD.n2198 AVDD.n2197 0.00970384
R4246 AVDD.n615 AVDD.n148 0.00967621
R4247 AVDD.n628 AVDD.n627 0.00947673
R4248 AVDD.n636 AVDD.n635 0.00947673
R4249 AVDD.n665 AVDD.n662 0.00947673
R4250 AVDD.n1475 AVDD.n1474 0.00947673
R4251 AVDD.n1370 AVDD.n1369 0.00947673
R4252 AVDD.n1362 AVDD.n1361 0.00947673
R4253 AVDD.n1334 AVDD.n1333 0.00947673
R4254 AVDD.n1326 AVDD.n1325 0.00947673
R4255 AVDD.n1117 AVDD.n958 0.00944828
R4256 AVDD.n649 AVDD.n648 0.00927724
R4257 AVDD.n650 AVDD.n649 0.00927724
R4258 AVDD.n1350 AVDD.n1349 0.00927724
R4259 AVDD.n1349 AVDD.n1345 0.00927724
R4260 AVDD.n630 AVDD.n142 0.00887828
R4261 AVDD.n1479 AVDD.n122 0.00887828
R4262 AVDD.n1367 AVDD.n1366 0.00887828
R4263 AVDD.n1331 AVDD.n1330 0.00887828
R4264 AVDD.n991 AVDD.n990 0.00877586
R4265 AVDD.n1178 AVDD.n744 0.00791176
R4266 AVDD.n1131 AVDD.n1130 0.00787705
R4267 AVDD.n992 AVDD.n991 0.00763793
R4268 AVDD.n396 AVDD.n395 0.00746812
R4269 AVDD.n521 AVDD.n513 0.00746812
R4270 AVDD.n942 AVDD.n941 0.0073513
R4271 AVDD.n784 AVDD.n783 0.0073513
R4272 AVDD.n755 AVDD.n754 0.0073513
R4273 AVDD.n948 AVDD.n756 0.0073513
R4274 AVDD.n947 AVDD.n946 0.0073513
R4275 AVDD.n760 AVDD.n758 0.0073513
R4276 AVDD.n779 AVDD.n778 0.0073513
R4277 AVDD.n775 AVDD.n764 0.0073513
R4278 AVDD.n774 AVDD.n773 0.0073513
R4279 AVDD.n772 AVDD.n765 0.0073513
R4280 AVDD.n945 AVDD.n781 0.00713029
R4281 AVDD.n761 AVDD.n757 0.00713029
R4282 AVDD.n939 AVDD.n785 0.0070075
R4283 AVDD.n938 AVDD.n782 0.0070075
R4284 AVDD.n768 AVDD.n767 0.0070075
R4285 AVDD.n770 AVDD.n769 0.0070075
R4286 AVDD.n1001 AVDD.n1000 0.00696552
R4287 AVDD.n921 AVDD.n920 0.00693383
R4288 AVDD.n924 AVDD.n906 0.00693383
R4289 AVDD.n927 AVDD.n925 0.00693383
R4290 AVDD.n926 AVDD.n904 0.00693383
R4291 AVDD.n929 AVDD.n928 0.00693383
R4292 AVDD.n808 AVDD.n801 0.00682401
R4293 AVDD.n1299 AVDD.n1247 0.00682401
R4294 AVDD.n762 AVDD.n759 0.00656548
R4295 AVDD.n952 AVDD.n753 0.00651637
R4296 AVDD.n1118 AVDD.n1117 0.0065
R4297 AVDD.n905 AVDD.n903 0.0064427
R4298 AVDD.n1314 AVDD.n1313 0.0063515
R4299 AVDD.n615 AVDD.n614 0.00598578
R4300 AVDD.n934 AVDD.n932 0.00595157
R4301 AVDD.n933 AVDD.n786 0.00595157
R4302 AVDD.n936 AVDD.n935 0.00595157
R4303 AVDD.n1226 AVDD.n714 0.00595157
R4304 AVDD.n1229 AVDD.n713 0.00595157
R4305 AVDD.n1002 AVDD.n1001 0.00531034
R4306 AVDD.n1082 AVDD.n1081 0.00512451
R4307 AVDD.n402 AVDD.n401 0.00509184
R4308 AVDD.n609 AVDD.n407 0.00509184
R4309 AVDD.n916 AVDD.n716 0.00489563
R4310 AVDD.n1004 AVDD.n1003 0.00484483
R4311 AVDD.n614 AVDD.n147 0.00445641
R4312 AVDD.n1950 AVDD.n59 0.00441304
R4313 AVDD.n1539 AVDD.n86 0.00441304
R4314 AVDD.n45 AVDD.n43 0.00441304
R4315 AVDD.n72 AVDD.n70 0.00441304
R4316 AVDD.n1936 AVDD.n1935 0.00429447
R4317 AVDD.n1525 AVDD.n1524 0.00429447
R4318 AVDD.n1745 AVDD.n1744 0.00429447
R4319 AVDD.n172 AVDD.n171 0.00429447
R4320 AVDD.n435 AVDD.n434 0.00418286
R4321 AVDD.n584 AVDD.n583 0.00418286
R4322 AVDD.n2182 AVDD.n19 0.00418286
R4323 AVDD.n1313 AVDD.n704 0.00409069
R4324 AVDD.n1028 AVDD.n1005 0.00355172
R4325 AVDD.n1224 AVDD.n1223 0.00342224
R4326 AVDD.n569 AVDD.n568 0.00334483
R4327 AVDD.n1225 AVDD.n1224 0.00302933
R4328 AVDD.n1067 AVDD.n992 0.00277586
R4329 AVDD.n1483 AVDD.n87 0.00272414
R4330 AVDD.n2140 AVDD.n2139 0.00272414
R4331 AVDD.n1032 AVDD.n1031 0.00267241
R4332 AVDD.n922 AVDD.n716 0.0025382
R4333 AVDD.n2178 AVDD.n2177 0.00237378
R4334 AVDD.n476 AVDD.n475 0.00237378
R4335 AVDD.n1404 AVDD.n118 0.00237378
R4336 AVDD.n1520 AVDD.n1519 0.00237378
R4337 AVDD.n508 AVDD.n506 0.00237378
R4338 AVDD.n825 AVDD.n824 0.00237378
R4339 AVDD.n846 AVDD.n844 0.00237378
R4340 AVDD.n1255 AVDD.n1253 0.00237378
R4341 AVDD.n1067 AVDD.n1066 0.00236207
R4342 AVDD.n2197 AVDD.n2196 0.0021987
R4343 AVDD.n925 AVDD.n924 0.00209618
R4344 AVDD.n934 AVDD.n933 0.00202251
R4345 AVDD.n936 AVDD.n786 0.00202251
R4346 AVDD.n935 AVDD.n785 0.00202251
R4347 AVDD.n769 AVDD.n714 0.00202251
R4348 AVDD.n1226 AVDD.n1225 0.00202251
R4349 AVDD.n1223 AVDD.n713 0.00202251
R4350 AVDD.n1032 AVDD.n752 0.00189655
R4351 AVDD.n1729 AVDD.n1728 0.00182807
R4352 AVDD.n1120 AVDD.n1119 0.00168966
R4353 AVDD.n2099 AVDD.n2098 0.00168421
R4354 AVDD.n2093 AVDD.n2092 0.00168421
R4355 AVDD.n2087 AVDD.n2086 0.00168421
R4356 AVDD.n2081 AVDD.n2080 0.00168421
R4357 AVDD.n1978 AVDD.n1977 0.00168421
R4358 AVDD.n1972 AVDD.n1971 0.00168421
R4359 AVDD.n1966 AVDD.n1965 0.00168421
R4360 AVDD.n2037 AVDD.n2036 0.00168421
R4361 AVDD.n2031 AVDD.n2030 0.00168421
R4362 AVDD.n2025 AVDD.n2024 0.00168421
R4363 AVDD.n2019 AVDD.n2018 0.00168421
R4364 AVDD.n2001 AVDD.n2000 0.00168421
R4365 AVDD.n1995 AVDD.n1994 0.00168421
R4366 AVDD.n1989 AVDD.n1988 0.00168421
R4367 AVDD.n1780 AVDD.n1776 0.00168421
R4368 AVDD.n1791 AVDD.n1789 0.00168421
R4369 AVDD.n1794 AVDD.n1785 0.00168421
R4370 AVDD.n1772 AVDD.n1768 0.00168421
R4371 AVDD.n1858 AVDD.n1765 0.00168421
R4372 AVDD.n1861 AVDD.n1761 0.00168421
R4373 AVDD.n1678 AVDD.n1580 0.00168421
R4374 AVDD.n1681 AVDD.n1576 0.00168421
R4375 AVDD.n1684 AVDD.n1572 0.00168421
R4376 AVDD.n1687 AVDD.n1568 0.00168421
R4377 AVDD.n1563 AVDD.n1562 0.00168421
R4378 AVDD.n1557 AVDD.n1556 0.00168421
R4379 AVDD.n1551 AVDD.n1550 0.00168421
R4380 AVDD.n1628 AVDD.n1627 0.00168421
R4381 AVDD.n1631 AVDD.n1623 0.00168421
R4382 AVDD.n1634 AVDD.n1619 0.00168421
R4383 AVDD.n1637 AVDD.n1615 0.00168421
R4384 AVDD.n1610 AVDD.n1609 0.00168421
R4385 AVDD.n1604 AVDD.n1603 0.00168421
R4386 AVDD.n1598 AVDD.n1597 0.00168421
R4387 AVDD.n230 AVDD.n226 0.00168421
R4388 AVDD.n222 AVDD.n221 0.00168421
R4389 AVDD.n216 AVDD.n215 0.00168421
R4390 AVDD.n287 AVDD.n283 0.00168421
R4391 AVDD.n279 AVDD.n278 0.00168421
R4392 AVDD.n273 AVDD.n272 0.00168421
R4393 AVDD.n1183 AVDD.n740 0.00168421
R4394 AVDD.n1186 AVDD.n736 0.00168421
R4395 AVDD.n1189 AVDD.n732 0.00168421
R4396 AVDD.n1192 AVDD.n728 0.00168421
R4397 AVDD.n1195 AVDD.n725 0.00168421
R4398 AVDD.n1198 AVDD.n721 0.00168421
R4399 AVDD.n1176 AVDD.n1173 0.00168421
R4400 AVDD.n1168 AVDD.n1165 0.00168421
R4401 AVDD.n1160 AVDD.n1157 0.00168421
R4402 AVDD.n1152 AVDD.n1150 0.00168421
R4403 AVDD.n1146 AVDD.n1143 0.00168421
R4404 AVDD.n1138 AVDD.n1135 0.00168421
R4405 AVDD.n1100 AVDD.n981 0.00168421
R4406 AVDD.n1103 AVDD.n977 0.00168421
R4407 AVDD.n1106 AVDD.n973 0.00168421
R4408 AVDD.n1109 AVDD.n969 0.00168421
R4409 AVDD.n1112 AVDD.n966 0.00168421
R4410 AVDD.n1115 AVDD.n962 0.00168421
R4411 AVDD.n142 AVDD.n140 0.00156391
R4412 AVDD.n1479 AVDD.n1478 0.00156391
R4413 AVDD.n1366 AVDD.n1365 0.00156391
R4414 AVDD.n1330 AVDD.n1329 0.00156391
R4415 AVDD.n1121 AVDD.n957 0.00153448
R4416 AVDD.n932 AVDD.n903 0.00153138
R4417 AVDD.n952 AVDD.n951 0.00133493
R4418 AVDD.n763 AVDD.n762 0.00128581
R4419 AVDD.n1030 AVDD.n1029 0.00106897
R4420 AVDD.n917 AVDD.n916 0.00104025
R4421 AVDD.n922 AVDD.n921 0.00104025
R4422 AVDD.n920 AVDD.n906 0.00104025
R4423 AVDD.n927 AVDD.n926 0.00104025
R4424 AVDD.n929 AVDD.n904 0.00104025
R4425 AVDD.n928 AVDD.n905 0.00104025
R4426 AVDD.n939 AVDD.n938 0.000966576
R4427 AVDD.n770 AVDD.n768 0.000966576
R4428 AVDD.n1057 AVDD.n1055 0.000762697
R4429 AVDD.n781 AVDD.n757 0.00072101
R4430 AVDD.n942 AVDD.n782 0.000622783
R4431 AVDD.n941 AVDD.n784 0.000622783
R4432 AVDD.n783 AVDD.n753 0.000622783
R4433 AVDD.n951 AVDD.n754 0.000622783
R4434 AVDD.n756 AVDD.n755 0.000622783
R4435 AVDD.n948 AVDD.n947 0.000622783
R4436 AVDD.n946 AVDD.n945 0.000622783
R4437 AVDD.n761 AVDD.n760 0.000622783
R4438 AVDD.n779 AVDD.n758 0.000622783
R4439 AVDD.n778 AVDD.n759 0.000622783
R4440 AVDD.n764 AVDD.n763 0.000622783
R4441 AVDD.n775 AVDD.n774 0.000622783
R4442 AVDD.n773 AVDD.n772 0.000622783
R4443 AVDD.n767 AVDD.n765 0.000622783
R4444 AVSS.n189 AVSS.n188 4252.69
R4445 AVSS.n473 AVSS.n472 661.869
R4446 AVSS.n429 AVSS.n192 661.869
R4447 AVSS.n426 AVSS.n74 661.869
R4448 AVSS.n76 AVSS.n75 656.895
R4449 AVSS.n469 AVSS.n190 656.895
R4450 AVSS.n476 AVSS.n73 656.895
R4451 AVSS.n472 AVSS.n76 656.434
R4452 AVSS.n469 AVSS.n192 656.434
R4453 AVSS.n476 AVSS.n74 656.434
R4454 AVSS.n473 AVSS.n75 653.672
R4455 AVSS.n429 AVSS.n190 653.672
R4456 AVSS.n426 AVSS.n73 653.672
R4457 AVSS.t34 AVSS.t82 517.433
R4458 AVSS.t49 AVSS.t138 517.433
R4459 AVSS.t99 AVSS.t4 454.447
R4460 AVSS.t31 AVSS.t178 450.327
R4461 AVSS.n124 AVSS.n91 383.618
R4462 AVSS.n164 AVSS.n91 381.962
R4463 AVSS.n124 AVSS.n90 381.132
R4464 AVSS.n164 AVSS.n90 379.474
R4465 AVSS.t133 AVSS.t34 329.651
R4466 AVSS.t138 AVSS.t96 329.651
R4467 AVSS.n124 AVSS.t49 275.635
R4468 AVSS.n188 AVSS.t4 275.495
R4469 AVSS.n166 AVSS.t31 275.495
R4470 AVSS.n165 AVSS.t82 275.495
R4471 AVSS.n167 AVSS.n79 267.474
R4472 AVSS.n187 AVSS.n79 266.829
R4473 AVSS.n167 AVSS.n78 266.276
R4474 AVSS.n187 AVSS.n78 265.632
R4475 AVSS.t96 AVSS.n123 244.294
R4476 AVSS.n123 AVSS.t133 233.7
R4477 AVSS.t235 AVSS.t77 178.191
R4478 AVSS.t172 AVSS.t46 178.191
R4479 AVSS.t144 AVSS.t201 173.123
R4480 AVSS.t19 AVSS.t175 173.123
R4481 AVSS.t178 AVSS.n89 168.946
R4482 AVSS.n89 AVSS.t99 160.706
R4483 AVSS.t58 AVSS.t158 158.528
R4484 AVSS.t67 AVSS.t28 158.528
R4485 AVSS.t2 AVSS.t114 155.487
R4486 AVSS.t13 AVSS.t25 155.487
R4487 AVSS.t10 AVSS.t235 113.523
R4488 AVSS.t201 AVSS.t10 113.523
R4489 AVSS.t222 AVSS.t144 113.523
R4490 AVSS.t175 AVSS.t43 113.523
R4491 AVSS.t43 AVSS.t172 113.523
R4492 AVSS.n470 AVSS.t19 109.469
R4493 AVSS.t16 AVSS.t163 95.8869
R4494 AVSS.t0 AVSS.t85 95.8869
R4495 AVSS.t77 AVSS.n426 94.9497
R4496 AVSS.t46 AVSS.n189 94.8732
R4497 AVSS.t70 AVSS.t22 93.8597
R4498 AVSS.t7 AVSS.t155 93.8597
R4499 AVSS.t37 AVSS.t55 90.8189
R4500 AVSS.n191 AVSS.t52 89.6025
R4501 AVSS.n166 AVSS.n165 84.7678
R4502 AVSS.n428 AVSS.t141 80.2775
R4503 AVSS.n475 AVSS.t1 80.2775
R4504 AVSS.n428 AVSS.n427 32.0302
R4505 AVSS.n475 AVSS.n474 29.1921
R4506 AVSS.t52 AVSS.t2 22.7051
R4507 AVSS.t25 AVSS.t37 22.7051
R4508 AVSS.t158 AVSS.t70 19.6643
R4509 AVSS.t22 AVSS.t7 19.6643
R4510 AVSS.t155 AVSS.t67 19.6643
R4511 AVSS.t114 AVSS.t16 17.6371
R4512 AVSS.t163 AVSS.t0 17.6371
R4513 AVSS.t85 AVSS.t13 17.6371
R4514 AVSS.t141 AVSS.t58 14.5963
R4515 AVSS.t28 AVSS.t1 14.5963
R4516 AVSS.n173 AVSS.t118 8.52542
R4517 AVSS.n92 AVSS.t81 8.52542
R4518 AVSS.n128 AVSS.t182 8.52542
R4519 AVSS.n132 AVSS.t213 8.52542
R4520 AVSS.n107 AVSS.t137 8.52542
R4521 AVSS.n115 AVSS.t95 8.52542
R4522 AVSS.n108 AVSS.t132 8.52542
R4523 AVSS.n109 AVSS.t211 8.52542
R4524 AVSS.n120 AVSS.t245 8.52542
R4525 AVSS.n122 AVSS.t203 8.52542
R4526 AVSS.n154 AVSS.t48 8.52542
R4527 AVSS.n152 AVSS.t74 8.52542
R4528 AVSS.n126 AVSS.t247 8.52542
R4529 AVSS.n147 AVSS.t180 8.52542
R4530 AVSS.n127 AVSS.t241 8.52542
R4531 AVSS.n141 AVSS.t33 8.52542
R4532 AVSS.n528 AVSS.t148 8.06917
R4533 AVSS.n239 AVSS.t12 8.06917
R4534 AVSS.n231 AVSS.t103 8.06917
R4535 AVSS.n229 AVSS.t15 8.06917
R4536 AVSS.n250 AVSS.t87 8.06917
R4537 AVSS.n224 AVSS.t165 8.06917
R4538 AVSS.n218 AVSS.t89 8.06917
R4539 AVSS.n261 AVSS.t66 8.06917
R4540 AVSS.n214 AVSS.t146 8.06917
R4541 AVSS.n212 AVSS.t69 8.06917
R4542 AVSS.n209 AVSS.t251 8.06917
R4543 AVSS.n2 AVSS.t54 8.06917
R4544 AVSS.n233 AVSS.t263 8.06917
R4545 AVSS.n240 AVSS.t84 8.06917
R4546 AVSS.n230 AVSS.t162 8.06917
R4547 AVSS.n228 AVSS.t113 8.06917
R4548 AVSS.n251 AVSS.t167 8.06917
R4549 AVSS.n217 AVSS.t79 8.06917
R4550 AVSS.n262 AVSS.t154 8.06917
R4551 AVSS.n213 AVSS.t259 8.06917
R4552 AVSS.n211 AVSS.t157 8.06917
R4553 AVSS.n208 AVSS.t140 8.06917
R4554 AVSS.n221 AVSS.t51 8.06917
R4555 AVSS.n220 AVSS.t111 8.06917
R4556 AVSS.n479 AVSS.t275 8.06917
R4557 AVSS.n480 AVSS.t126 8.06917
R4558 AVSS.n482 AVSS.t215 8.06917
R4559 AVSS.n221 AVSS.t230 8.06917
R4560 AVSS.n220 AVSS.t271 8.06917
R4561 AVSS.n479 AVSS.t184 8.06917
R4562 AVSS.n480 AVSS.t27 8.06917
R4563 AVSS.n482 AVSS.t116 8.06917
R4564 AVSS.n297 AVSS.t205 8.06917
R4565 AVSS.n301 AVSS.t21 8.06917
R4566 AVSS.n296 AVSS.t207 8.06917
R4567 AVSS.n295 AVSS.t188 8.06917
R4568 AVSS.n309 AVSS.t257 8.06917
R4569 AVSS.n294 AVSS.t190 8.06917
R4570 AVSS.n293 AVSS.t243 8.06917
R4571 AVSS.n316 AVSS.t72 8.06917
R4572 AVSS.n292 AVSS.t267 8.06917
R4573 AVSS.n386 AVSS.t224 8.06917
R4574 AVSS.n389 AVSS.t42 8.06917
R4575 AVSS.n385 AVSS.t226 8.06917
R4576 AVSS.n394 AVSS.t18 8.06917
R4577 AVSS.n397 AVSS.t105 8.06917
R4578 AVSS.n384 AVSS.t24 8.06917
R4579 AVSS.n383 AVSS.t120 8.06917
R4580 AVSS.n404 AVSS.t209 8.06917
R4581 AVSS.n382 AVSS.t130 8.06917
R4582 AVSS.n9 AVSS.t124 8.06917
R4583 AVSS.n512 AVSS.t93 8.06917
R4584 AVSS.n5 AVSS.t171 8.06917
R4585 AVSS.n517 AVSS.t269 8.06917
R4586 AVSS.n4 AVSS.t174 8.06917
R4587 AVSS.n522 AVSS.t261 8.06917
R4588 AVSS.n6 AVSS.t237 8.06917
R4589 AVSS.n6 AVSS.t281 8.06917
R4590 AVSS.n6 AVSS.t194 8.06917
R4591 AVSS.n6 AVSS.t45 8.06917
R4592 AVSS.n435 AVSS.t122 8.06917
R4593 AVSS.n433 AVSS.t273 8.06917
R4594 AVSS.n432 AVSS.t135 8.06917
R4595 AVSS.n204 AVSS.t57 8.06917
R4596 AVSS.n205 AVSS.t160 8.06917
R4597 AVSS.n193 AVSS.t150 8.06917
R4598 AVSS.n455 AVSS.t232 8.06917
R4599 AVSS.n194 AVSS.t152 8.06917
R4600 AVSS.n195 AVSS.t217 8.06917
R4601 AVSS.n447 AVSS.t39 8.06917
R4602 AVSS.n196 AVSS.t219 8.06917
R4603 AVSS.n197 AVSS.t196 8.06917
R4604 AVSS.n440 AVSS.t6 8.06917
R4605 AVSS.n198 AVSS.t198 8.06917
R4606 AVSS.n460 AVSS.t36 8.06917
R4607 AVSS.n462 AVSS.t192 8.06917
R4608 AVSS.n463 AVSS.t62 8.06917
R4609 AVSS.n466 AVSS.t239 8.06917
R4610 AVSS.n465 AVSS.t91 8.06917
R4611 AVSS.n275 AVSS.t221 8.06917
R4612 AVSS.n202 AVSS.t143 8.06917
R4613 AVSS.n201 AVSS.t200 8.06917
R4614 AVSS.n282 AVSS.t9 8.06917
R4615 AVSS.n200 AVSS.t234 8.06917
R4616 AVSS.n287 AVSS.t128 8.06917
R4617 AVSS.n289 AVSS.t279 8.06917
R4618 AVSS.n290 AVSS.t76 8.06917
R4619 AVSS.n423 AVSS.t249 8.06917
R4620 AVSS.n422 AVSS.t107 8.06917
R4621 AVSS.n420 AVSS.t169 8.06917
R4622 AVSS.n342 AVSS.t324 6.72766
R4623 AVSS.n81 AVSS.t3 6.60917
R4624 AVSS.n81 AVSS.t253 6.60917
R4625 AVSS.n81 AVSS.t64 6.60917
R4626 AVSS.n81 AVSS.t101 6.60917
R4627 AVSS.n81 AVSS.t277 6.60917
R4628 AVSS.n179 AVSS.t186 6.60917
R4629 AVSS.n85 AVSS.t109 6.60917
R4630 AVSS.n133 AVSS.t177 6.60917
R4631 AVSS.n84 AVSS.t98 6.60917
R4632 AVSS.n174 AVSS.t265 6.60917
R4633 AVSS.n171 AVSS.t228 6.60917
R4634 AVSS.n88 AVSS.t30 6.60917
R4635 AVSS.n93 AVSS.t60 6.60917
R4636 AVSS.n129 AVSS.t255 6.60917
R4637 AVSS.n38 AVSS.n35 6.53862
R4638 AVSS.n83 AVSS.n82 5.49372
R4639 AVSS.n339 AVSS.t374 5.47432
R4640 AVSS.n333 AVSS.n332 5.31981
R4641 AVSS.n43 AVSS.t307 5.28484
R4642 AVSS.n51 AVSS.n50 5.28484
R4643 AVSS.n42 AVSS.t284 5.28484
R4644 AVSS.n338 AVSS.n320 5.26136
R4645 AVSS.t5 AVSS.n184 5.2505
R4646 AVSS.n185 AVSS.t5 5.2505
R4647 AVSS.n184 AVSS.t254 5.2505
R4648 AVSS.n185 AVSS.t254 5.2505
R4649 AVSS.n184 AVSS.t65 5.2505
R4650 AVSS.n185 AVSS.t65 5.2505
R4651 AVSS.n184 AVSS.t102 5.2505
R4652 AVSS.n185 AVSS.t102 5.2505
R4653 AVSS.n184 AVSS.t278 5.2505
R4654 AVSS.n185 AVSS.t278 5.2505
R4655 AVSS.n178 AVSS.t187 5.2505
R4656 AVSS.n182 AVSS.t110 5.2505
R4657 AVSS.t100 AVSS.n83 5.2505
R4658 AVSS.n137 AVSS.t179 5.2505
R4659 AVSS.n68 AVSS.n67 5.16888
R4660 AVSS.n21 AVSS.n20 5.15456
R4661 AVSS.n411 AVSS.n410 5.09675
R4662 AVSS.n501 AVSS.n497 4.63106
R4663 AVSS.n491 AVSS.n487 4.63106
R4664 AVSS.n29 AVSS.n25 4.63106
R4665 AVSS.n334 AVSS.n333 4.61712
R4666 AVSS.n415 AVSS.n414 4.61712
R4667 AVSS.n158 AVSS.n157 4.61585
R4668 AVSS.n161 AVSS.n160 4.61585
R4669 AVSS.n413 AVSS.n412 4.61078
R4670 AVSS.n505 AVSS.n503 4.61078
R4671 AVSS.n495 AVSS.n493 4.61078
R4672 AVSS.n33 AVSS.n31 4.61078
R4673 AVSS.n23 AVSS.n21 4.61078
R4674 AVSS.n412 AVSS.n411 4.60825
R4675 AVSS.n506 AVSS.n505 4.60825
R4676 AVSS.n496 AVSS.n495 4.60825
R4677 AVSS.n34 AVSS.n33 4.60825
R4678 AVSS.n24 AVSS.n23 4.60825
R4679 AVSS.n343 AVSS.n339 4.60439
R4680 AVSS.n157 AVSS.n156 4.60318
R4681 AVSS.n160 AVSS.n159 4.60318
R4682 AVSS.n335 AVSS.n334 4.60191
R4683 AVSS.n416 AVSS.n415 4.60191
R4684 AVSS.n502 AVSS.n501 4.58796
R4685 AVSS.n492 AVSS.n491 4.58796
R4686 AVSS.n30 AVSS.n29 4.58796
R4687 AVSS.n323 AVSS.n321 4.5005
R4688 AVSS.n327 AVSS.n324 4.5005
R4689 AVSS.n330 AVSS.n328 4.5005
R4690 AVSS.n22 AVSS.n18 4.5005
R4691 AVSS.n28 AVSS.n17 4.5005
R4692 AVSS.n32 AVSS.n16 4.5005
R4693 AVSS.n490 AVSS.n15 4.5005
R4694 AVSS.n494 AVSS.n14 4.5005
R4695 AVSS.n500 AVSS.n13 4.5005
R4696 AVSS.n504 AVSS.n12 4.5005
R4697 AVSS.n98 AVSS.n95 4.5005
R4698 AVSS.n104 AVSS.n101 4.5005
R4699 AVSS.n362 AVSS.t339 4.41563
R4700 AVSS.n377 AVSS.n375 4.41563
R4701 AVSS.n360 AVSS.t290 4.41563
R4702 AVSS.n346 AVSS.n344 4.41563
R4703 AVSS.n60 AVSS.t305 4.22616
R4704 AVSS.n58 AVSS.t337 4.22616
R4705 AVSS.n342 AVSS.n341 4.21432
R4706 AVSS.n338 AVSS.n337 4.21432
R4707 AVSS.n474 AVSS.t40 4.05489
R4708 AVSS.n46 AVSS.n45 4.02484
R4709 AVSS.n49 AVSS.n48 4.02484
R4710 AVSS.n41 AVSS.n40 4.02484
R4711 AVSS.n38 AVSS.n37 4.02484
R4712 AVSS.n60 AVSS.t333 4.02247
R4713 AVSS.n58 AVSS.t388 4.02247
R4714 AVSS.n330 AVSS.n329 4.00471
R4715 AVSS.n323 AVSS.n322 4.00471
R4716 AVSS.n61 AVSS.n11 3.96014
R4717 AVSS.n362 AVSS.t306 3.833
R4718 AVSS.n377 AVSS.n376 3.833
R4719 AVSS.n360 AVSS.t384 3.833
R4720 AVSS.n346 AVSS.n345 3.833
R4721 AVSS.n504 AVSS.t377 3.81405
R4722 AVSS.n494 AVSS.t375 3.81405
R4723 AVSS.n32 AVSS.t381 3.81405
R4724 AVSS.n22 AVSS.t370 3.81405
R4725 AVSS.n359 AVSS.n353 3.80578
R4726 AVSS.n374 AVSS.n368 3.80578
R4727 AVSS.n41 AVSS.n38 3.80578
R4728 AVSS.n49 AVSS.n46 3.80578
R4729 AVSS.n417 AVSS.n416 3.76738
R4730 AVSS.n510 AVSS.t125 3.37683
R4731 AVSS.t149 AVSS.n1 3.3605
R4732 AVSS.n234 AVSS.t149 3.3605
R4733 AVSS.n236 AVSS.t14 3.3605
R4734 AVSS.t17 AVSS.n227 3.3605
R4735 AVSS.n248 AVSS.t88 3.3605
R4736 AVSS.t90 AVSS.n216 3.3605
R4737 AVSS.n258 AVSS.t68 3.3605
R4738 AVSS.t71 AVSS.n210 3.3605
R4739 AVSS.n270 AVSS.t252 3.3605
R4740 AVSS.t252 AVSS.n203 3.3605
R4741 AVSS.n235 AVSS.t264 3.3605
R4742 AVSS.n238 AVSS.t86 3.3605
R4743 AVSS.n247 AVSS.t115 3.3605
R4744 AVSS.n249 AVSS.t168 3.3605
R4745 AVSS.t168 AVSS.n226 3.3605
R4746 AVSS.t80 AVSS.n256 3.3605
R4747 AVSS.n257 AVSS.t80 3.3605
R4748 AVSS.n260 AVSS.t156 3.3605
R4749 AVSS.n269 AVSS.t159 3.3605
R4750 AVSS.t142 AVSS.n271 3.3605
R4751 AVSS.t206 AVSS.n298 3.3605
R4752 AVSS.n304 AVSS.t208 3.3605
R4753 AVSS.t189 AVSS.n305 3.3605
R4754 AVSS.n312 AVSS.t191 3.3605
R4755 AVSS.t244 AVSS.n313 3.3605
R4756 AVSS.n319 AVSS.t268 3.3605
R4757 AVSS.t225 AVSS.n10 3.3605
R4758 AVSS.n392 AVSS.t227 3.3605
R4759 AVSS.n393 AVSS.t20 3.3605
R4760 AVSS.n400 AVSS.t26 3.3605
R4761 AVSS.t121 AVSS.n401 3.3605
R4762 AVSS.n407 AVSS.t131 3.3605
R4763 AVSS.t125 AVSS.n509 3.3605
R4764 AVSS.t173 AVSS.n514 3.3605
R4765 AVSS.n520 AVSS.t176 3.3605
R4766 AVSS.n521 AVSS.t262 3.3605
R4767 AVSS.n8 AVSS.t282 3.3605
R4768 AVSS.t282 AVSS.n7 3.3605
R4769 AVSS.n8 AVSS.t195 3.3605
R4770 AVSS.n7 AVSS.t195 3.3605
R4771 AVSS.n8 AVSS.t47 3.3605
R4772 AVSS.n7 AVSS.t47 3.3605
R4773 AVSS.n458 AVSS.t151 3.3605
R4774 AVSS.t153 AVSS.n452 3.3605
R4775 AVSS.n451 AVSS.t218 3.3605
R4776 AVSS.t220 AVSS.n444 3.3605
R4777 AVSS.n443 AVSS.t197 3.3605
R4778 AVSS.t199 AVSS.n437 3.3605
R4779 AVSS.n278 AVSS.t145 3.3605
R4780 AVSS.t202 AVSS.n279 3.3605
R4781 AVSS.n285 AVSS.t236 3.3605
R4782 AVSS.n367 AVSS.n364 3.15563
R4783 AVSS.n373 AVSS.n370 3.15563
R4784 AVSS.n358 AVSS.n355 3.15563
R4785 AVSS.n352 AVSS.n349 3.15563
R4786 AVSS.n136 AVSS.n135 3.1505
R4787 AVSS.n181 AVSS.n180 3.1505
R4788 AVSS.n343 AVSS.n342 3.02463
R4789 AVSS.n66 AVSS.n63 2.96616
R4790 AVSS.n57 AVSS.n54 2.96616
R4791 AVSS.n25 AVSS.n24 2.885
R4792 AVSS.n497 AVSS.n496 2.885
R4793 AVSS.n471 AVSS.n470 2.83857
R4794 AVSS.n487 AVSS.n486 2.795
R4795 AVSS.n66 AVSS.n65 2.76247
R4796 AVSS.n57 AVSS.n56 2.76247
R4797 AVSS.n327 AVSS.n326 2.74471
R4798 AVSS.n59 AVSS.n57 2.71914
R4799 AVSS.n368 AVSS.n362 2.71872
R4800 AVSS.n118 AVSS.t139 2.6955
R4801 AVSS.n114 AVSS.t97 2.6955
R4802 AVSS.n112 AVSS.t134 2.6955
R4803 AVSS.t212 AVSS.n87 2.6955
R4804 AVSS.n150 AVSS.t248 2.6955
R4805 AVSS.n146 AVSS.t181 2.6955
R4806 AVSS.n144 AVSS.t242 2.6955
R4807 AVSS.n140 AVSS.t35 2.6955
R4808 AVSS.n177 AVSS.t266 2.6255
R4809 AVSS.n172 AVSS.t229 2.6255
R4810 AVSS.n170 AVSS.t32 2.6255
R4811 AVSS.n94 AVSS.t61 2.6255
R4812 AVSS.n131 AVSS.t256 2.6255
R4813 AVSS.n367 AVSS.n366 2.573
R4814 AVSS.n373 AVSS.n372 2.573
R4815 AVSS.n358 AVSS.n357 2.573
R4816 AVSS.n352 AVSS.n351 2.573
R4817 AVSS.n500 AVSS.n499 2.55405
R4818 AVSS.n490 AVSS.n489 2.55405
R4819 AVSS.n28 AVSS.n27 2.55405
R4820 AVSS.n68 AVSS.n59 2.46014
R4821 AVSS.n162 AVSS.n161 2.45973
R4822 AVSS.n156 AVSS.n155 2.45073
R4823 AVSS.n379 AVSS.n361 2.38034
R4824 AVSS.n43 AVSS.n11 2.37491
R4825 AVSS.n52 AVSS.n51 2.32143
R4826 AVSS.n484 AVSS.n483 2.30076
R4827 AVSS.n410 AVSS.n335 2.26738
R4828 AVSS.n380 AVSS.n343 2.23722
R4829 AVSS.n104 AVSS.n103 2.15932
R4830 AVSS.n98 AVSS.n97 2.15932
R4831 AVSS.n157 AVSS.n106 2.15458
R4832 AVSS.n160 AVSS.n100 2.15458
R4833 AVSS.n69 AVSS.n52 2.13932
R4834 AVSS.n524 AVSS.n523 2.1005
R4835 AVSS.n519 AVSS.n518 2.1005
R4836 AVSS.n516 AVSS.n515 2.1005
R4837 AVSS.t110 AVSS.n181 2.1005
R4838 AVSS.n181 AVSS.t187 2.1005
R4839 AVSS.n136 AVSS.t100 2.1005
R4840 AVSS.t179 AVSS.n136 2.1005
R4841 AVSS.n439 AVSS.n438 2.1005
R4842 AVSS.n442 AVSS.n441 2.1005
R4843 AVSS.n446 AVSS.n445 2.1005
R4844 AVSS.n450 AVSS.n449 2.1005
R4845 AVSS.n454 AVSS.n453 2.1005
R4846 AVSS.n457 AVSS.n456 2.1005
R4847 AVSS.n284 AVSS.n283 2.1005
R4848 AVSS.n281 AVSS.n280 2.1005
R4849 AVSS.n277 AVSS.n276 2.1005
R4850 AVSS.n406 AVSS.n405 2.1005
R4851 AVSS.n403 AVSS.n402 2.1005
R4852 AVSS.n399 AVSS.n398 2.1005
R4853 AVSS.n396 AVSS.n395 2.1005
R4854 AVSS.n391 AVSS.n390 2.1005
R4855 AVSS.n388 AVSS.n387 2.1005
R4856 AVSS.n318 AVSS.n317 2.1005
R4857 AVSS.n315 AVSS.n314 2.1005
R4858 AVSS.n311 AVSS.n310 2.1005
R4859 AVSS.n307 AVSS.n306 2.1005
R4860 AVSS.n303 AVSS.n302 2.1005
R4861 AVSS.n300 AVSS.n299 2.1005
R4862 AVSS.n273 AVSS.n272 2.1005
R4863 AVSS.n268 AVSS.n267 2.1005
R4864 AVSS.n259 AVSS.n215 2.1005
R4865 AVSS.n246 AVSS.n245 2.1005
R4866 AVSS.n237 AVSS.n232 2.1005
R4867 AVSS.n526 AVSS.n525 2.1005
R4868 AVSS.n266 AVSS.n265 2.1005
R4869 AVSS.n264 AVSS.n263 2.1005
R4870 AVSS.n255 AVSS.n254 2.1005
R4871 AVSS.n253 AVSS.n252 2.1005
R4872 AVSS.n244 AVSS.n243 2.1005
R4873 AVSS.n242 AVSS.n241 2.1005
R4874 AVSS.n508 AVSS.n507 1.7274
R4875 AVSS.n222 AVSS.t53 1.6805
R4876 AVSS.n219 AVSS.t112 1.6805
R4877 AVSS.n478 AVSS.t276 1.6805
R4878 AVSS.n481 AVSS.t127 1.6805
R4879 AVSS.n71 AVSS.t216 1.6805
R4880 AVSS.n222 AVSS.t231 1.6805
R4881 AVSS.n219 AVSS.t272 1.6805
R4882 AVSS.n478 AVSS.t185 1.6805
R4883 AVSS.n481 AVSS.t29 1.6805
R4884 AVSS.n71 AVSS.t117 1.6805
R4885 AVSS.n513 AVSS.t94 1.6805
R4886 AVSS.n511 AVSS.t238 1.6805
R4887 AVSS.n436 AVSS.t123 1.6805
R4888 AVSS.n434 AVSS.t274 1.6805
R4889 AVSS.n431 AVSS.t136 1.6805
R4890 AVSS.n199 AVSS.t59 1.6805
R4891 AVSS.n206 AVSS.t161 1.6805
R4892 AVSS.n459 AVSS.t38 1.6805
R4893 AVSS.n461 AVSS.t193 1.6805
R4894 AVSS.n464 AVSS.t63 1.6805
R4895 AVSS.n467 AVSS.t240 1.6805
R4896 AVSS.n0 AVSS.t92 1.6805
R4897 AVSS.n286 AVSS.t129 1.6805
R4898 AVSS.n288 AVSS.t280 1.6805
R4899 AVSS.n291 AVSS.t78 1.6805
R4900 AVSS.n424 AVSS.t250 1.6805
R4901 AVSS.n421 AVSS.t108 1.6805
R4902 AVSS.n419 AVSS.t170 1.6805
R4903 AVSS.n418 AVSS.n417 1.67828
R4904 AVSS.n409 AVSS.n408 1.67828
R4905 AVSS.n347 AVSS.n320 1.67718
R4906 AVSS.n507 AVSS.n506 1.60175
R4907 AVSS.n143 AVSS.n142 1.5755
R4908 AVSS.n149 AVSS.n148 1.5755
R4909 AVSS.n111 AVSS.n110 1.5755
R4910 AVSS.n117 AVSS.n116 1.5755
R4911 AVSS.n410 AVSS.n409 1.5005
R4912 AVSS.n380 AVSS.n379 1.5005
R4913 AVSS.n486 AVSS.n485 1.5005
R4914 AVSS.n69 AVSS.n68 1.5005
R4915 AVSS.n61 AVSS.n60 1.46537
R4916 AVSS.n67 AVSS.n66 1.46537
R4917 AVSS.n59 AVSS.n58 1.46537
R4918 AVSS.n368 AVSS.n367 1.46537
R4919 AVSS.n374 AVSS.n373 1.46537
R4920 AVSS.n378 AVSS.n377 1.46537
R4921 AVSS.n361 AVSS.n360 1.46537
R4922 AVSS.n359 AVSS.n358 1.46537
R4923 AVSS.n353 AVSS.n352 1.46537
R4924 AVSS.n347 AVSS.n346 1.46537
R4925 AVSS.n175 AVSS.t119 1.348
R4926 AVSS.n169 AVSS.t83 1.348
R4927 AVSS.n130 AVSS.t183 1.348
R4928 AVSS.n139 AVSS.t214 1.348
R4929 AVSS.n119 AVSS.t246 1.348
R4930 AVSS.n121 AVSS.t204 1.348
R4931 AVSS.n153 AVSS.t50 1.348
R4932 AVSS.n151 AVSS.t75 1.348
R4933 AVSS.n159 AVSS.n158 1.265
R4934 AVSS.t104 AVSS.n242 1.2605
R4935 AVSS.n242 AVSS.t14 1.2605
R4936 AVSS.n243 AVSS.t17 1.2605
R4937 AVSS.n243 AVSS.t104 1.2605
R4938 AVSS.t166 AVSS.n253 1.2605
R4939 AVSS.n253 AVSS.t88 1.2605
R4940 AVSS.n254 AVSS.t90 1.2605
R4941 AVSS.n254 AVSS.t166 1.2605
R4942 AVSS.t147 AVSS.n264 1.2605
R4943 AVSS.n264 AVSS.t68 1.2605
R4944 AVSS.n265 AVSS.t71 1.2605
R4945 AVSS.n265 AVSS.t147 1.2605
R4946 AVSS.n525 AVSS.t264 1.2605
R4947 AVSS.n525 AVSS.t56 1.2605
R4948 AVSS.n237 AVSS.t164 1.2605
R4949 AVSS.t86 AVSS.n237 1.2605
R4950 AVSS.t115 AVSS.n246 1.2605
R4951 AVSS.n246 AVSS.t164 1.2605
R4952 AVSS.n259 AVSS.t260 1.2605
R4953 AVSS.t156 AVSS.n259 1.2605
R4954 AVSS.t159 AVSS.n268 1.2605
R4955 AVSS.n268 AVSS.t260 1.2605
R4956 AVSS.n272 AVSS.t223 1.2605
R4957 AVSS.n272 AVSS.t142 1.2605
R4958 AVSS.n299 AVSS.t23 1.2605
R4959 AVSS.n299 AVSS.t206 1.2605
R4960 AVSS.t208 AVSS.n303 1.2605
R4961 AVSS.n303 AVSS.t23 1.2605
R4962 AVSS.n306 AVSS.t258 1.2605
R4963 AVSS.n306 AVSS.t189 1.2605
R4964 AVSS.t191 AVSS.n311 1.2605
R4965 AVSS.n311 AVSS.t258 1.2605
R4966 AVSS.n314 AVSS.t73 1.2605
R4967 AVSS.n314 AVSS.t244 1.2605
R4968 AVSS.t268 AVSS.n318 1.2605
R4969 AVSS.n318 AVSS.t73 1.2605
R4970 AVSS.n387 AVSS.t44 1.2605
R4971 AVSS.n387 AVSS.t225 1.2605
R4972 AVSS.t227 AVSS.n391 1.2605
R4973 AVSS.n391 AVSS.t44 1.2605
R4974 AVSS.t106 AVSS.n396 1.2605
R4975 AVSS.n396 AVSS.t20 1.2605
R4976 AVSS.t26 AVSS.n399 1.2605
R4977 AVSS.n399 AVSS.t106 1.2605
R4978 AVSS.n402 AVSS.t210 1.2605
R4979 AVSS.n402 AVSS.t121 1.2605
R4980 AVSS.t131 AVSS.n406 1.2605
R4981 AVSS.n406 AVSS.t210 1.2605
R4982 AVSS.n332 AVSS.t385 1.2605
R4983 AVSS.n332 AVSS.n331 1.2605
R4984 AVSS.n326 AVSS.t365 1.2605
R4985 AVSS.n326 AVSS.n325 1.2605
R4986 AVSS.n364 AVSS.t338 1.2605
R4987 AVSS.n364 AVSS.n363 1.2605
R4988 AVSS.n366 AVSS.t376 1.2605
R4989 AVSS.n366 AVSS.n365 1.2605
R4990 AVSS.n370 AVSS.t318 1.2605
R4991 AVSS.n370 AVSS.n369 1.2605
R4992 AVSS.n372 AVSS.t397 1.2605
R4993 AVSS.n372 AVSS.n371 1.2605
R4994 AVSS.n355 AVSS.t289 1.2605
R4995 AVSS.n355 AVSS.n354 1.2605
R4996 AVSS.n357 AVSS.t398 1.2605
R4997 AVSS.n357 AVSS.n356 1.2605
R4998 AVSS.n349 AVSS.t350 1.2605
R4999 AVSS.n349 AVSS.n348 1.2605
R5000 AVSS.n351 AVSS.t298 1.2605
R5001 AVSS.n351 AVSS.n350 1.2605
R5002 AVSS.n341 AVSS.t323 1.2605
R5003 AVSS.n341 AVSS.n340 1.2605
R5004 AVSS.n337 AVSS.t373 1.2605
R5005 AVSS.n337 AVSS.n336 1.2605
R5006 AVSS.n63 AVSS.t304 1.2605
R5007 AVSS.n63 AVSS.n62 1.2605
R5008 AVSS.n65 AVSS.t291 1.2605
R5009 AVSS.n65 AVSS.n64 1.2605
R5010 AVSS.n54 AVSS.t336 1.2605
R5011 AVSS.n54 AVSS.n53 1.2605
R5012 AVSS.n56 AVSS.t387 1.2605
R5013 AVSS.n56 AVSS.n55 1.2605
R5014 AVSS.n45 AVSS.t364 1.2605
R5015 AVSS.n45 AVSS.n44 1.2605
R5016 AVSS.n48 AVSS.t311 1.2605
R5017 AVSS.n48 AVSS.n47 1.2605
R5018 AVSS.n40 AVSS.t283 1.2605
R5019 AVSS.n40 AVSS.n39 1.2605
R5020 AVSS.n37 AVSS.t349 1.2605
R5021 AVSS.n37 AVSS.n36 1.2605
R5022 AVSS.n499 AVSS.t299 1.2605
R5023 AVSS.n499 AVSS.n498 1.2605
R5024 AVSS.n489 AVSS.t363 1.2605
R5025 AVSS.n489 AVSS.n488 1.2605
R5026 AVSS.n27 AVSS.t380 1.2605
R5027 AVSS.n27 AVSS.n26 1.2605
R5028 AVSS.n20 AVSS.t346 1.2605
R5029 AVSS.n20 AVSS.n19 1.2605
R5030 AVSS.n515 AVSS.t270 1.2605
R5031 AVSS.n515 AVSS.t173 1.2605
R5032 AVSS.t176 AVSS.n519 1.2605
R5033 AVSS.n519 AVSS.t270 1.2605
R5034 AVSS.t56 AVSS.n524 1.2605
R5035 AVSS.n524 AVSS.t262 1.2605
R5036 AVSS.n457 AVSS.t233 1.2605
R5037 AVSS.t151 AVSS.n457 1.2605
R5038 AVSS.n453 AVSS.t153 1.2605
R5039 AVSS.n453 AVSS.t233 1.2605
R5040 AVSS.n450 AVSS.t41 1.2605
R5041 AVSS.t218 AVSS.n450 1.2605
R5042 AVSS.n445 AVSS.t220 1.2605
R5043 AVSS.n445 AVSS.t41 1.2605
R5044 AVSS.n442 AVSS.t8 1.2605
R5045 AVSS.t197 AVSS.n442 1.2605
R5046 AVSS.n438 AVSS.t199 1.2605
R5047 AVSS.n438 AVSS.t8 1.2605
R5048 AVSS.t145 AVSS.n277 1.2605
R5049 AVSS.n277 AVSS.t223 1.2605
R5050 AVSS.n280 AVSS.t11 1.2605
R5051 AVSS.n280 AVSS.t202 1.2605
R5052 AVSS.t236 AVSS.n284 1.2605
R5053 AVSS.n284 AVSS.t11 1.2605
R5054 AVSS.n353 AVSS.n347 1.25428
R5055 AVSS.n361 AVSS.n359 1.25428
R5056 AVSS.n378 AVSS.n374 1.25428
R5057 AVSS.n339 AVSS.n338 1.25428
R5058 AVSS.n42 AVSS.n41 1.25428
R5059 AVSS.n51 AVSS.n49 1.25428
R5060 AVSS.n46 AVSS.n43 1.25428
R5061 AVSS.n67 AVSS.n61 1.25428
R5062 AVSS.n427 AVSS.t222 1.21682
R5063 AVSS.n191 AVSS.t40 1.21682
R5064 AVSS.n471 AVSS.t55 1.21682
R5065 AVSS.n484 AVSS.n70 1.13691
R5066 AVSS.n117 AVSS.t97 1.1205
R5067 AVSS.t139 AVSS.n117 1.1205
R5068 AVSS.n111 AVSS.t212 1.1205
R5069 AVSS.t134 AVSS.n111 1.1205
R5070 AVSS.n103 AVSS.t310 1.1205
R5071 AVSS.n103 AVSS.n102 1.1205
R5072 AVSS.n106 AVSS.t371 1.1205
R5073 AVSS.n106 AVSS.n105 1.1205
R5074 AVSS.n97 AVSS.t372 1.1205
R5075 AVSS.n97 AVSS.n96 1.1205
R5076 AVSS.n100 AVSS.t386 1.1205
R5077 AVSS.n100 AVSS.n99 1.1205
R5078 AVSS.n149 AVSS.t181 1.1205
R5079 AVSS.t248 AVSS.n149 1.1205
R5080 AVSS.n143 AVSS.t35 1.1205
R5081 AVSS.t242 AVSS.n143 1.1205
R5082 AVSS.n31 AVSS.n30 0.9995
R5083 AVSS.n493 AVSS.n492 0.9995
R5084 AVSS.n503 AVSS.n502 0.9995
R5085 AVSS.n414 AVSS.n413 0.973625
R5086 AVSS.n485 AVSS.n484 0.970331
R5087 AVSS.n417 AVSS.n320 0.585196
R5088 AVSS.n409 AVSS.n380 0.585196
R5089 AVSS.n485 AVSS.n69 0.585196
R5090 AVSS.n507 AVSS.n11 0.585196
R5091 AVSS.n186 AVSS.n80 0.239651
R5092 AVSS.n52 AVSS.n42 0.236091
R5093 AVSS.n168 AVSS.n167 0.186214
R5094 AVSS.n167 AVSS.n166 0.186214
R5095 AVSS.n187 AVSS.n186 0.186214
R5096 AVSS.n188 AVSS.n187 0.186214
R5097 AVSS.n379 AVSS.n378 0.177184
R5098 AVSS.n134 AVSS.n79 0.163
R5099 AVSS.n89 AVSS.n79 0.163
R5100 AVSS.n86 AVSS.n78 0.163
R5101 AVSS.n89 AVSS.n78 0.163
R5102 AVSS.n125 AVSS.n124 0.141041
R5103 AVSS.n164 AVSS.n163 0.141041
R5104 AVSS.n165 AVSS.n164 0.141041
R5105 AVSS.n416 AVSS.n321 0.14
R5106 AVSS.n414 AVSS.n321 0.14
R5107 AVSS.n413 AVSS.n324 0.14
R5108 AVSS.n411 AVSS.n324 0.14
R5109 AVSS.n335 AVSS.n328 0.14
R5110 AVSS.n333 AVSS.n328 0.14
R5111 AVSS.n21 AVSS.n18 0.14
R5112 AVSS.n24 AVSS.n18 0.14
R5113 AVSS.n25 AVSS.n17 0.14
R5114 AVSS.n30 AVSS.n17 0.14
R5115 AVSS.n31 AVSS.n16 0.14
R5116 AVSS.n34 AVSS.n16 0.14
R5117 AVSS.n487 AVSS.n15 0.14
R5118 AVSS.n492 AVSS.n15 0.14
R5119 AVSS.n493 AVSS.n14 0.14
R5120 AVSS.n496 AVSS.n14 0.14
R5121 AVSS.n497 AVSS.n13 0.14
R5122 AVSS.n502 AVSS.n13 0.14
R5123 AVSS.n503 AVSS.n12 0.14
R5124 AVSS.n506 AVSS.n12 0.14
R5125 AVSS.n161 AVSS.n95 0.14
R5126 AVSS.n159 AVSS.n95 0.14
R5127 AVSS.n158 AVSS.n101 0.14
R5128 AVSS.n156 AVSS.n101 0.14
R5129 AVSS.n183 AVSS.n83 0.132207
R5130 AVSS.n145 AVSS.n91 0.108833
R5131 AVSS.n123 AVSS.n91 0.108833
R5132 AVSS.n113 AVSS.n90 0.108833
R5133 AVSS.n123 AVSS.n90 0.108833
R5134 AVSS.n512 AVSS.n511 0.105988
R5135 AVSS.n461 AVSS.n460 0.105988
R5136 AVSS.n435 AVSS.n434 0.105988
R5137 AVSS.n288 AVSS.n287 0.105988
R5138 AVSS.n421 AVSS.n420 0.105988
R5139 AVSS.n527 AVSS.n0 0.102012
R5140 AVSS.n207 AVSS.n206 0.102012
R5141 AVSS.n486 AVSS.n34 0.10175
R5142 AVSS.n183 AVSS.n84 0.100659
R5143 AVSS.n426 AVSS.n425 0.0769706
R5144 AVSS.n430 AVSS.n429 0.0769706
R5145 AVSS.n429 AVSS.n428 0.0769706
R5146 AVSS.n469 AVSS.n468 0.0769706
R5147 AVSS.n470 AVSS.n469 0.0769706
R5148 AVSS.n80 AVSS.n76 0.0769706
R5149 AVSS.n189 AVSS.n76 0.0769706
R5150 AVSS.n477 AVSS.n476 0.0769706
R5151 AVSS.n476 AVSS.n475 0.0769706
R5152 AVSS.n473 AVSS.n72 0.0769706
R5153 AVSS.n474 AVSS.n473 0.0769706
R5154 AVSS.n430 AVSS.n199 0.072814
R5155 AVSS.n425 AVSS.n424 0.072814
R5156 AVSS.n121 AVSS.n120 0.0718609
R5157 AVSS.n153 AVSS.n152 0.0718609
R5158 AVSS.n468 AVSS.n464 0.0681047
R5159 AVSS.n468 AVSS.n467 0.0678953
R5160 AVSS.n274 AVSS.n73 0.0646975
R5161 AVSS.n427 AVSS.n73 0.0646975
R5162 AVSS.n448 AVSS.n190 0.0646975
R5163 AVSS.n191 AVSS.n190 0.0646975
R5164 AVSS.n472 AVSS.n77 0.0646975
R5165 AVSS.n472 AVSS.n471 0.0646975
R5166 AVSS.n308 AVSS.n74 0.0646975
R5167 AVSS.n427 AVSS.n74 0.0646975
R5168 AVSS.n75 AVSS.n3 0.0646975
R5169 AVSS.n471 AVSS.n75 0.0646975
R5170 AVSS.n225 AVSS.n192 0.0646975
R5171 AVSS.n192 AVSS.n191 0.0646975
R5172 AVSS.n431 AVSS.n430 0.063186
R5173 AVSS.n425 AVSS.n291 0.063186
R5174 AVSS.n482 AVSS.n481 0.0533671
R5175 AVSS.n223 AVSS.n222 0.0513741
R5176 AVSS.n182 AVSS.n85 0.0431396
R5177 AVSS.n180 AVSS.n179 0.0431396
R5178 AVSS.n179 AVSS.n178 0.0431396
R5179 AVSS.n86 AVSS.n85 0.0420736
R5180 AVSS.n463 AVSS.n462 0.041314
R5181 AVSS.n433 AVSS.n432 0.041314
R5182 AVSS.n290 AVSS.n289 0.041314
R5183 AVSS.n466 AVSS.n465 0.0411047
R5184 AVSS.n205 AVSS.n204 0.0411047
R5185 AVSS.n423 AVSS.n422 0.0411047
R5186 AVSS.n514 AVSS.n513 0.039811
R5187 AVSS.n286 AVSS.n285 0.039811
R5188 AVSS.n459 AVSS.n458 0.0385295
R5189 AVSS.n437 AVSS.n436 0.0385295
R5190 AVSS.n151 AVSS.n150 0.0365464
R5191 AVSS.n119 AVSS.n118 0.0364399
R5192 AVSS.n401 AVSS.n400 0.0354077
R5193 AVSS.n393 AVSS.n392 0.0354077
R5194 AVSS.n313 AVSS.n312 0.0354077
R5195 AVSS.n305 AVSS.n304 0.0354077
R5196 AVSS.n444 AVSS.n443 0.0353617
R5197 AVSS.n452 AVSS.n451 0.0353617
R5198 AVSS.n120 AVSS.n119 0.0346894
R5199 AVSS.n122 AVSS.n121 0.0346894
R5200 AVSS.n154 AVSS.n153 0.0346894
R5201 AVSS.n152 AVSS.n151 0.0346894
R5202 AVSS.n478 AVSS.n477 0.0342762
R5203 AVSS.n140 AVSS.n139 0.0342758
R5204 AVSS.n407 AVSS.n382 0.0337454
R5205 AVSS.n405 AVSS.n382 0.0337454
R5206 AVSS.n405 AVSS.n404 0.0337454
R5207 AVSS.n404 AVSS.n403 0.0337454
R5208 AVSS.n403 AVSS.n383 0.0337454
R5209 AVSS.n401 AVSS.n383 0.0337454
R5210 AVSS.n400 AVSS.n384 0.0337454
R5211 AVSS.n398 AVSS.n384 0.0337454
R5212 AVSS.n398 AVSS.n397 0.0337454
R5213 AVSS.n395 AVSS.n394 0.0337454
R5214 AVSS.n394 AVSS.n393 0.0337454
R5215 AVSS.n392 AVSS.n385 0.0337454
R5216 AVSS.n390 AVSS.n385 0.0337454
R5217 AVSS.n390 AVSS.n389 0.0337454
R5218 AVSS.n389 AVSS.n388 0.0337454
R5219 AVSS.n388 AVSS.n386 0.0337454
R5220 AVSS.n386 AVSS.n10 0.0337454
R5221 AVSS.n319 AVSS.n292 0.0337454
R5222 AVSS.n317 AVSS.n292 0.0337454
R5223 AVSS.n317 AVSS.n316 0.0337454
R5224 AVSS.n316 AVSS.n315 0.0337454
R5225 AVSS.n315 AVSS.n293 0.0337454
R5226 AVSS.n313 AVSS.n293 0.0337454
R5227 AVSS.n312 AVSS.n294 0.0337454
R5228 AVSS.n310 AVSS.n294 0.0337454
R5229 AVSS.n310 AVSS.n309 0.0337454
R5230 AVSS.n307 AVSS.n295 0.0337454
R5231 AVSS.n305 AVSS.n295 0.0337454
R5232 AVSS.n304 AVSS.n296 0.0337454
R5233 AVSS.n302 AVSS.n296 0.0337454
R5234 AVSS.n302 AVSS.n301 0.0337454
R5235 AVSS.n301 AVSS.n300 0.0337454
R5236 AVSS.n300 AVSS.n297 0.0337454
R5237 AVSS.n298 AVSS.n297 0.0337454
R5238 AVSS.n437 AVSS.n198 0.0337016
R5239 AVSS.n439 AVSS.n198 0.0337016
R5240 AVSS.n440 AVSS.n439 0.0337016
R5241 AVSS.n441 AVSS.n440 0.0337016
R5242 AVSS.n441 AVSS.n197 0.0337016
R5243 AVSS.n443 AVSS.n197 0.0337016
R5244 AVSS.n444 AVSS.n196 0.0337016
R5245 AVSS.n446 AVSS.n196 0.0337016
R5246 AVSS.n447 AVSS.n446 0.0337016
R5247 AVSS.n449 AVSS.n195 0.0337016
R5248 AVSS.n451 AVSS.n195 0.0337016
R5249 AVSS.n452 AVSS.n194 0.0337016
R5250 AVSS.n454 AVSS.n194 0.0337016
R5251 AVSS.n455 AVSS.n454 0.0337016
R5252 AVSS.n456 AVSS.n455 0.0337016
R5253 AVSS.n456 AVSS.n193 0.0337016
R5254 AVSS.n458 AVSS.n193 0.0337016
R5255 AVSS.n395 AVSS.n77 0.033033
R5256 AVSS.n308 AVSS.n307 0.033033
R5257 AVSS.n449 AVSS.n448 0.0329901
R5258 AVSS.n176 AVSS.n87 0.032073
R5259 AVSS.n141 AVSS.n140 0.0319607
R5260 AVSS.n142 AVSS.n141 0.0319607
R5261 AVSS.n142 AVSS.n127 0.0319607
R5262 AVSS.n144 AVSS.n127 0.0319607
R5263 AVSS.n147 AVSS.n146 0.0319607
R5264 AVSS.n148 AVSS.n147 0.0319607
R5265 AVSS.n148 AVSS.n126 0.0319607
R5266 AVSS.n150 AVSS.n126 0.0319607
R5267 AVSS.n109 AVSS.n87 0.0319607
R5268 AVSS.n110 AVSS.n109 0.0319607
R5269 AVSS.n110 AVSS.n108 0.0319607
R5270 AVSS.n112 AVSS.n108 0.0319607
R5271 AVSS.n115 AVSS.n114 0.0319607
R5272 AVSS.n116 AVSS.n115 0.0319607
R5273 AVSS.n116 AVSS.n107 0.0319607
R5274 AVSS.n118 AVSS.n107 0.0319607
R5275 AVSS.n219 AVSS.n72 0.0319161
R5276 AVSS.n521 AVSS.n520 0.0315563
R5277 AVSS.n279 AVSS.n278 0.0315563
R5278 AVSS.n513 AVSS.n512 0.0314767
R5279 AVSS.n460 AVSS.n459 0.0314767
R5280 AVSS.n462 AVSS.n461 0.0314767
R5281 AVSS.n464 AVSS.n463 0.0314767
R5282 AVSS.n467 AVSS.n466 0.0314767
R5283 AVSS.n465 AVSS.n0 0.0314767
R5284 AVSS.n436 AVSS.n435 0.0314767
R5285 AVSS.n434 AVSS.n433 0.0314767
R5286 AVSS.n432 AVSS.n431 0.0314767
R5287 AVSS.n204 AVSS.n199 0.0314767
R5288 AVSS.n206 AVSS.n205 0.0314767
R5289 AVSS.n287 AVSS.n286 0.0314767
R5290 AVSS.n289 AVSS.n288 0.0314767
R5291 AVSS.n291 AVSS.n290 0.0314767
R5292 AVSS.n424 AVSS.n423 0.0314767
R5293 AVSS.n422 AVSS.n421 0.0314767
R5294 AVSS.n420 AVSS.n419 0.0314767
R5295 AVSS.n523 AVSS.n522 0.0300775
R5296 AVSS.n522 AVSS.n521 0.0300775
R5297 AVSS.n520 AVSS.n4 0.0300775
R5298 AVSS.n518 AVSS.n4 0.0300775
R5299 AVSS.n518 AVSS.n517 0.0300775
R5300 AVSS.n517 AVSS.n516 0.0300775
R5301 AVSS.n516 AVSS.n5 0.0300775
R5302 AVSS.n514 AVSS.n5 0.0300775
R5303 AVSS.n285 AVSS.n200 0.0300775
R5304 AVSS.n283 AVSS.n200 0.0300775
R5305 AVSS.n283 AVSS.n282 0.0300775
R5306 AVSS.n282 AVSS.n281 0.0300775
R5307 AVSS.n281 AVSS.n201 0.0300775
R5308 AVSS.n279 AVSS.n201 0.0300775
R5309 AVSS.n278 AVSS.n202 0.0300775
R5310 AVSS.n276 AVSS.n202 0.0300775
R5311 AVSS.n276 AVSS.n275 0.0300775
R5312 AVSS.n178 AVSS.n177 0.0280818
R5313 AVSS.n509 AVSS.n9 0.0277138
R5314 AVSS.n508 AVSS.n10 0.0271502
R5315 AVSS.n183 AVSS.n182 0.0259315
R5316 AVSS.n132 AVSS.n131 0.0255699
R5317 AVSS.n523 AVSS.n3 0.0231186
R5318 AVSS.n511 AVSS.n510 0.0217442
R5319 AVSS.n419 AVSS.n418 0.0213083
R5320 AVSS.n221 AVSS.n220 0.0209545
R5321 AVSS.n480 AVSS.n479 0.0208496
R5322 AVSS.n408 AVSS.n407 0.0206172
R5323 AVSS.n418 AVSS.n319 0.0206172
R5324 AVSS.n298 AVSS.n70 0.0204409
R5325 AVSS.n155 AVSS.n154 0.0185
R5326 AVSS.n171 AVSS.n170 0.0181748
R5327 AVSS.n135 AVSS.n133 0.0173337
R5328 AVSS.n137 AVSS.n133 0.0173337
R5329 AVSS.n125 AVSS.n122 0.0172219
R5330 AVSS.n134 AVSS.n84 0.0169128
R5331 AVSS.n408 AVSS.n381 0.016599
R5332 AVSS.n139 AVSS.n138 0.0164441
R5333 AVSS.n129 AVSS.n128 0.0160769
R5334 AVSS.n222 AVSS.n221 0.0160245
R5335 AVSS.n220 AVSS.n219 0.0160245
R5336 AVSS.n479 AVSS.n478 0.0160245
R5337 AVSS.n481 AVSS.n480 0.0160245
R5338 AVSS.n381 AVSS.n70 0.0158871
R5339 AVSS.n274 AVSS.n273 0.0157873
R5340 AVSS.n146 AVSS.n145 0.0156685
R5341 AVSS.n114 AVSS.n113 0.0156685
R5342 AVSS.n509 AVSS.n508 0.0137679
R5343 AVSS.n145 AVSS.n144 0.0136461
R5344 AVSS.n113 AVSS.n112 0.0136461
R5345 AVSS.n172 AVSS.n171 0.0118287
R5346 AVSS.n174 AVSS.n173 0.011514
R5347 AVSS.n510 AVSS.n9 0.0113855
R5348 AVSS.n483 AVSS.n71 0.0113305
R5349 AVSS.n131 AVSS.n130 0.0105699
R5350 AVSS.n138 AVSS.n137 0.0105401
R5351 AVSS.n168 AVSS.n88 0.00999301
R5352 AVSS.n270 AVSS.n269 0.00799437
R5353 AVSS.n258 AVSS.n257 0.00799437
R5354 AVSS.n271 AVSS.n209 0.00752176
R5355 AVSS.n217 AVSS.n216 0.00752176
R5356 AVSS.n256 AVSS.n218 0.00752176
R5357 AVSS.n248 AVSS.n247 0.007488
R5358 AVSS.n236 AVSS.n235 0.007488
R5359 AVSS.n162 AVSS.n94 0.00721329
R5360 AVSS.n7 AVSS.n6 0.00704376
R5361 AVSS.n185 AVSS.n81 0.00704376
R5362 AVSS.n184 AVSS.n81 0.00704376
R5363 AVSS.n228 AVSS.n227 0.00701538
R5364 AVSS.n245 AVSS.n229 0.00701538
R5365 AVSS.n244 AVSS.n230 0.00701538
R5366 AVSS.n232 AVSS.n231 0.00701538
R5367 AVSS.n241 AVSS.n240 0.00701538
R5368 AVSS.n239 AVSS.n238 0.00701538
R5369 AVSS.n255 AVSS.n223 0.00684659
R5370 AVSS.n211 AVSS.n210 0.00667779
R5371 AVSS.n267 AVSS.n212 0.00667779
R5372 AVSS.n266 AVSS.n213 0.00667779
R5373 AVSS.n215 AVSS.n214 0.00667779
R5374 AVSS.n263 AVSS.n262 0.00667779
R5375 AVSS.n261 AVSS.n260 0.00667779
R5376 AVSS.n173 AVSS.n172 0.00653147
R5377 AVSS.n175 AVSS.n174 0.00632168
R5378 AVSS.n483 AVSS.n482 0.00619059
R5379 AVSS.n207 AVSS.n203 0.00617142
R5380 AVSS.n252 AVSS.n251 0.00617142
R5381 AVSS.n250 AVSS.n249 0.00617142
R5382 AVSS.n234 AVSS.n233 0.00617142
R5383 AVSS.n2 AVSS.n1 0.00617142
R5384 AVSS.n92 AVSS.n88 0.00611189
R5385 AVSS.n226 AVSS.n225 0.00596887
R5386 AVSS.n93 AVSS.n92 0.00490559
R5387 AVSS.n80 AVSS.n8 0.00489366
R5388 AVSS.n186 AVSS.n185 0.00489366
R5389 AVSS.n510 AVSS.n8 0.00442625
R5390 AVSS.n163 AVSS.n93 0.00432867
R5391 AVSS.n252 AVSS.n226 0.00428095
R5392 AVSS.n251 AVSS.n250 0.00428095
R5393 AVSS.n249 AVSS.n248 0.00428095
R5394 AVSS.n235 AVSS.n234 0.00428095
R5395 AVSS.n528 AVSS.n527 0.00428095
R5396 AVSS.n526 AVSS.n1 0.00428095
R5397 AVSS.n177 AVSS.n176 0.00385664
R5398 AVSS.n269 AVSS.n210 0.00377457
R5399 AVSS.n212 AVSS.n211 0.00377457
R5400 AVSS.n267 AVSS.n266 0.00377457
R5401 AVSS.n214 AVSS.n213 0.00377457
R5402 AVSS.n263 AVSS.n215 0.00377457
R5403 AVSS.n262 AVSS.n261 0.00377457
R5404 AVSS.n260 AVSS.n258 0.00377457
R5405 AVSS.n233 AVSS 0.00370705
R5406 AVSS.n224 AVSS.n223 0.00360578
R5407 AVSS.n247 AVSS.n227 0.00343698
R5408 AVSS.n229 AVSS.n228 0.00343698
R5409 AVSS.n245 AVSS.n244 0.00343698
R5410 AVSS.n231 AVSS.n230 0.00343698
R5411 AVSS.n241 AVSS.n232 0.00343698
R5412 AVSS.n240 AVSS.n239 0.00343698
R5413 AVSS.n238 AVSS.n236 0.00343698
R5414 AVSS.n510 AVSS.n6 0.0031175
R5415 AVSS.n477 AVSS.n72 0.00296504
R5416 AVSS.n273 AVSS.n203 0.00293061
R5417 AVSS.n209 AVSS.n208 0.00293061
R5418 AVSS.n271 AVSS.n270 0.00293061
R5419 AVSS.n257 AVSS.n216 0.00293061
R5420 AVSS.n218 AVSS.n217 0.00293061
R5421 AVSS.n256 AVSS.n255 0.00293061
R5422 AVSS.n381 AVSS.n71 0.00286014
R5423 AVSS.n176 AVSS.n175 0.00265035
R5424 AVSS.n128 AVSS.n94 0.00265035
R5425 AVSS.n527 AVSS.n526 0.00239047
R5426 AVSS.n169 AVSS.n168 0.00223077
R5427 AVSS.n155 AVSS.n125 0.00209763
R5428 AVSS.n208 AVSS.n207 0.00185034
R5429 AVSS.n130 AVSS.n129 0.00175874
R5430 AVSS.n334 AVSS.n330 0.00168421
R5431 AVSS.n412 AVSS.n327 0.00168421
R5432 AVSS.n415 AVSS.n323 0.00168421
R5433 AVSS.n505 AVSS.n504 0.00168421
R5434 AVSS.n501 AVSS.n500 0.00168421
R5435 AVSS.n495 AVSS.n494 0.00168421
R5436 AVSS.n491 AVSS.n490 0.00168421
R5437 AVSS.n33 AVSS.n32 0.00168421
R5438 AVSS.n29 AVSS.n28 0.00168421
R5439 AVSS.n23 AVSS.n22 0.00168421
R5440 AVSS.n157 AVSS.n104 0.00168421
R5441 AVSS.n160 AVSS.n98 0.00168421
R5442 AVSS.n180 AVSS.n86 0.00156599
R5443 AVSS.n184 AVSS.n183 0.00155167
R5444 AVSS.n138 AVSS.n132 0.00139161
R5445 AVSS.n163 AVSS.n162 0.00128671
R5446 AVSS.n397 AVSS.n77 0.0012124
R5447 AVSS.n309 AVSS.n308 0.0012124
R5448 AVSS.n448 AVSS.n447 0.00121146
R5449 AVSS.n275 AVSS.n274 0.0011338
R5450 AVSS.n528 AVSS 0.00107389
R5451 AVSS.n135 AVSS.n134 0.000920842
R5452 AVSS.n225 AVSS.n224 0.000702551
R5453 AVSS.n3 AVSS.n2 0.000702551
R5454 AVSS.n170 AVSS.n169 0.000604895
R5455 a_5396_n6451.n380 a_5396_n6451.t260 8.38704
R5456 a_5396_n6451.n374 a_5396_n6451.t255 8.38704
R5457 a_5396_n6451.n168 a_5396_n6451.t195 8.46135
R5458 a_5396_n6451.n170 a_5396_n6451.t123 8.46135
R5459 a_5396_n6451.n43 a_5396_n6451.t127 8.48081
R5460 a_5396_n6451.n38 a_5396_n6451.t173 8.48081
R5461 a_5396_n6451.n21 a_5396_n6451.t179 8.10567
R5462 a_5396_n6451.n26 a_5396_n6451.t111 8.10567
R5463 a_5396_n6451.n26 a_5396_n6451.t203 8.10567
R5464 a_5396_n6451.n223 a_5396_n6451.t197 8.10567
R5465 a_5396_n6451.n248 a_5396_n6451.t250 8.10567
R5466 a_5396_n6451.n203 a_5396_n6451.t108 8.10567
R5467 a_5396_n6451.n204 a_5396_n6451.t275 8.10567
R5468 a_5396_n6451.n227 a_5396_n6451.t149 8.10567
R5469 a_5396_n6451.n226 a_5396_n6451.t139 8.10567
R5470 a_5396_n6451.n207 a_5396_n6451.t191 8.10567
R5471 a_5396_n6451.n208 a_5396_n6451.t245 8.10567
R5472 a_5396_n6451.n230 a_5396_n6451.t233 8.10567
R5473 a_5396_n6451.n253 a_5396_n6451.t110 8.10567
R5474 a_5396_n6451.n28 a_5396_n6451.t166 8.10567
R5475 a_5396_n6451.n28 a_5396_n6451.t157 8.10567
R5476 a_5396_n6451.n288 a_5396_n6451.t208 8.10567
R5477 a_5396_n6451.n30 a_5396_n6451.t251 8.10567
R5478 a_5396_n6451.n30 a_5396_n6451.t239 8.10567
R5479 a_5396_n6451.n200 a_5396_n6451.t118 8.10567
R5480 a_5396_n6451.n21 a_5396_n6451.t171 8.10567
R5481 a_5396_n6451.n211 a_5396_n6451.t248 8.10567
R5482 a_5396_n6451.n234 a_5396_n6451.t235 8.10567
R5483 a_5396_n6451.n278 a_5396_n6451.t237 8.10567
R5484 a_5396_n6451.n171 a_5396_n6451.t209 8.10567
R5485 a_5396_n6451.n171 a_5396_n6451.t270 8.10567
R5486 a_5396_n6451.n3 a_5396_n6451.t229 8.10567
R5487 a_5396_n6451.n3 a_5396_n6451.t172 8.10567
R5488 a_5396_n6451.n173 a_5396_n6451.t257 8.10567
R5489 a_5396_n6451.n174 a_5396_n6451.t214 8.10567
R5490 a_5396_n6451.n0 a_5396_n6451.t142 8.10567
R5491 a_5396_n6451.n0 a_5396_n6451.t279 8.10567
R5492 a_5396_n6451.n281 a_5396_n6451.t185 8.10567
R5493 a_5396_n6451.n177 a_5396_n6451.t129 8.10567
R5494 a_5396_n6451.n6 a_5396_n6451.t253 8.10567
R5495 a_5396_n6451.n6 a_5396_n6451.t188 8.10567
R5496 a_5396_n6451.n159 a_5396_n6451.t163 8.10567
R5497 a_5396_n6451.n159 a_5396_n6451.t126 8.10567
R5498 a_5396_n6451.n300 a_5396_n6451.t242 8.10567
R5499 a_5396_n6451.n161 a_5396_n6451.t136 8.10567
R5500 a_5396_n6451.n161 a_5396_n6451.t274 8.10567
R5501 a_5396_n6451.n286 a_5396_n6451.t216 8.10567
R5502 a_5396_n6451.n181 a_5396_n6451.t199 8.10567
R5503 a_5396_n6451.n180 a_5396_n6451.t158 8.10567
R5504 a_5396_n6451.n180 a_5396_n6451.t121 8.10567
R5505 a_5396_n6451.n18 a_5396_n6451.t226 8.10567
R5506 a_5396_n6451.n24 a_5396_n6451.t198 8.10567
R5507 a_5396_n6451.n24 a_5396_n6451.t261 8.10567
R5508 a_5396_n6451.n236 a_5396_n6451.t218 8.10567
R5509 a_5396_n6451.n256 a_5396_n6451.t161 8.10567
R5510 a_5396_n6451.n213 a_5396_n6451.t244 8.10567
R5511 a_5396_n6451.n214 a_5396_n6451.t204 8.10567
R5512 a_5396_n6451.n212 a_5396_n6451.t133 8.10567
R5513 a_5396_n6451.n239 a_5396_n6451.t271 8.10567
R5514 a_5396_n6451.n218 a_5396_n6451.t174 8.10567
R5515 a_5396_n6451.n219 a_5396_n6451.t119 8.10567
R5516 a_5396_n6451.n217 a_5396_n6451.t236 8.10567
R5517 a_5396_n6451.n242 a_5396_n6451.t181 8.10567
R5518 a_5396_n6451.n32 a_5396_n6451.t138 8.10567
R5519 a_5396_n6451.n32 a_5396_n6451.t278 8.10567
R5520 a_5396_n6451.n201 a_5396_n6451.t220 8.10567
R5521 a_5396_n6451.n34 a_5396_n6451.t117 8.10567
R5522 a_5396_n6451.n34 a_5396_n6451.t254 8.10567
R5523 a_5396_n6451.n202 a_5396_n6451.t193 8.10567
R5524 a_5396_n6451.n18 a_5396_n6451.t187 8.10567
R5525 a_5396_n6451.n222 a_5396_n6451.t147 8.10567
R5526 a_5396_n6451.n246 a_5396_n6451.t109 8.10567
R5527 a_5396_n6451.n194 a_5396_n6451.t165 8.10567
R5528 a_5396_n6451.n184 a_5396_n6451.t135 8.10567
R5529 a_5396_n6451.n184 a_5396_n6451.t196 8.10567
R5530 a_5396_n6451.n9 a_5396_n6451.t156 8.10567
R5531 a_5396_n6451.n9 a_5396_n6451.t273 8.10567
R5532 a_5396_n6451.n275 a_5396_n6451.t182 8.10567
R5533 a_5396_n6451.n186 a_5396_n6451.t145 8.10567
R5534 a_5396_n6451.n12 a_5396_n6451.t246 8.10567
R5535 a_5396_n6451.n12 a_5396_n6451.t205 8.10567
R5536 a_5396_n6451.n189 a_5396_n6451.t114 8.10567
R5537 a_5396_n6451.n190 a_5396_n6451.t228 8.10567
R5538 a_5396_n6451.n15 a_5396_n6451.t176 8.10567
R5539 a_5396_n6451.n15 a_5396_n6451.t120 8.10567
R5540 a_5396_n6451.n163 a_5396_n6451.t269 8.10567
R5541 a_5396_n6451.n163 a_5396_n6451.t225 8.10567
R5542 a_5396_n6451.n287 a_5396_n6451.t169 8.10567
R5543 a_5396_n6451.n165 a_5396_n6451.t240 8.10567
R5544 a_5396_n6451.n165 a_5396_n6451.t202 8.10567
R5545 a_5396_n6451.n304 a_5396_n6451.t146 8.10567
R5546 a_5396_n6451.n195 a_5396_n6451.t130 8.10567
R5547 a_5396_n6451.n193 a_5396_n6451.t264 8.10567
R5548 a_5396_n6451.n193 a_5396_n6451.t222 8.10567
R5549 a_5396_n6451.n89 a_5396_n6451.t124 8.10567
R5550 a_5396_n6451.n91 a_5396_n6451.t116 8.10567
R5551 a_5396_n6451.n94 a_5396_n6451.t164 8.10567
R5552 a_5396_n6451.n367 a_5396_n6451.t154 8.10567
R5553 a_5396_n6451.n479 a_5396_n6451.t151 8.10567
R5554 a_5396_n6451.n478 a_5396_n6451.t141 8.10567
R5555 a_5396_n6451.n477 a_5396_n6451.t192 8.10567
R5556 a_5396_n6451.n42 a_5396_n6451.t219 8.10567
R5557 a_5396_n6451.n98 a_5396_n6451.t210 8.10567
R5558 a_5396_n6451.n99 a_5396_n6451.t266 8.10567
R5559 a_5396_n6451.n71 a_5396_n6451.t194 8.10567
R5560 a_5396_n6451.n74 a_5396_n6451.t186 8.10567
R5561 a_5396_n6451.n373 a_5396_n6451.t265 8.10567
R5562 a_5396_n6451.n472 a_5396_n6451.t232 8.10567
R5563 a_5396_n6451.n471 a_5396_n6451.t224 8.10567
R5564 a_5396_n6451.n470 a_5396_n6451.t276 8.10567
R5565 a_5396_n6451.n40 a_5396_n6451.t207 8.10567
R5566 a_5396_n6451.n77 a_5396_n6451.t262 8.10567
R5567 a_5396_n6451.n80 a_5396_n6451.t252 8.10567
R5568 a_5396_n6451.n83 a_5396_n6451.t125 8.10567
R5569 a_5396_n6451.n115 a_5396_n6451.t238 8.10567
R5570 a_5396_n6451.n157 a_5396_n6451.t200 8.10567
R5571 a_5396_n6451.n140 a_5396_n6451.t128 8.10567
R5572 a_5396_n6451.n311 a_5396_n6451.t267 8.10567
R5573 a_5396_n6451.n410 a_5396_n6451.t178 8.10567
R5574 a_5396_n6451.n409 a_5396_n6451.t137 8.10567
R5575 a_5396_n6451.n408 a_5396_n6451.t259 8.10567
R5576 a_5396_n6451.n167 a_5396_n6451.t256 8.10567
R5577 a_5396_n6451.n142 a_5396_n6451.t213 8.10567
R5578 a_5396_n6451.n125 a_5396_n6451.t155 8.10567
R5579 a_5396_n6451.n109 a_5396_n6451.t223 8.10567
R5580 a_5396_n6451.n152 a_5396_n6451.t184 8.10567
R5581 a_5396_n6451.n306 a_5396_n6451.t144 8.10567
R5582 a_5396_n6451.n397 a_5396_n6451.t153 8.10567
R5583 a_5396_n6451.n396 a_5396_n6451.t115 8.10567
R5584 a_5396_n6451.n395 a_5396_n6451.t231 8.10567
R5585 a_5396_n6451.n317 a_5396_n6451.t170 8.10567
R5586 a_5396_n6451.n156 a_5396_n6451.t112 8.10567
R5587 a_5396_n6451.n136 a_5396_n6451.t234 8.10567
R5588 a_5396_n6451.n122 a_5396_n6451.t175 8.10567
R5589 a_5396_n6451.n60 a_5396_n6451.t215 8.10567
R5590 a_5396_n6451.n62 a_5396_n6451.t177 8.10567
R5591 a_5396_n6451.n64 a_5396_n6451.t106 8.10567
R5592 a_5396_n6451.n427 a_5396_n6451.t241 8.10567
R5593 a_5396_n6451.n419 a_5396_n6451.t168 8.10567
R5594 a_5396_n6451.n420 a_5396_n6451.t132 8.10567
R5595 a_5396_n6451.n421 a_5396_n6451.t249 8.10567
R5596 a_5396_n6451.n39 a_5396_n6451.t230 8.10567
R5597 a_5396_n6451.n66 a_5396_n6451.t190 8.10567
R5598 a_5396_n6451.n68 a_5396_n6451.t134 8.10567
R5599 a_5396_n6451.n48 a_5396_n6451.t201 8.10567
R5600 a_5396_n6451.n50 a_5396_n6451.t162 8.10567
R5601 a_5396_n6451.n379 a_5396_n6451.t122 8.10567
R5602 a_5396_n6451.n385 a_5396_n6451.t143 8.10567
R5603 a_5396_n6451.n384 a_5396_n6451.t280 8.10567
R5604 a_5396_n6451.n383 a_5396_n6451.t221 8.10567
R5605 a_5396_n6451.n36 a_5396_n6451.t148 8.10567
R5606 a_5396_n6451.n52 a_5396_n6451.t268 8.10567
R5607 a_5396_n6451.n57 a_5396_n6451.t211 8.10567
R5608 a_5396_n6451.n58 a_5396_n6451.t152 8.10567
R5609 a_5396_n6451.n106 a_5396_n6451.t167 8.10567
R5610 a_5396_n6451.n150 a_5396_n6451.t131 8.10567
R5611 a_5396_n6451.n131 a_5396_n6451.t227 8.10567
R5612 a_5396_n6451.n314 a_5396_n6451.t189 8.10567
R5613 a_5396_n6451.n447 a_5396_n6451.t107 8.10567
R5614 a_5396_n6451.n448 a_5396_n6451.t243 8.10567
R5615 a_5396_n6451.n449 a_5396_n6451.t183 8.10567
R5616 a_5396_n6451.n169 a_5396_n6451.t180 8.10567
R5617 a_5396_n6451.n134 a_5396_n6451.t140 8.10567
R5618 a_5396_n6451.n120 a_5396_n6451.t263 8.10567
R5619 a_5396_n6451.n105 a_5396_n6451.t150 8.10567
R5620 a_5396_n6451.n144 a_5396_n6451.t113 8.10567
R5621 a_5396_n6451.n310 a_5396_n6451.t247 8.10567
R5622 a_5396_n6451.n439 a_5396_n6451.t258 8.10567
R5623 a_5396_n6451.n438 a_5396_n6451.t217 8.10567
R5624 a_5396_n6451.n437 a_5396_n6451.t159 8.10567
R5625 a_5396_n6451.n319 a_5396_n6451.t272 8.10567
R5626 a_5396_n6451.n147 a_5396_n6451.t212 8.10567
R5627 a_5396_n6451.n128 a_5396_n6451.t160 8.10567
R5628 a_5396_n6451.n117 a_5396_n6451.t277 8.10567
R5629 a_5396_n6451.n575 a_5396_n6451.n571 7.22198
R5630 a_5396_n6451.n613 a_5396_n6451.n349 7.22198
R5631 a_5396_n6451.n488 a_5396_n6451.n485 6.77653
R5632 a_5396_n6451.n586 a_5396_n6451.n583 6.77653
R5633 a_5396_n6451.n507 a_5396_n6451.t30 6.7761
R5634 a_5396_n6451.n605 a_5396_n6451.t13 6.7761
R5635 a_5396_n6451.n341 a_5396_n6451.n527 6.86989
R5636 a_5396_n6451.n330 a_5396_n6451.n352 6.77231
R5637 a_5396_n6451.n340 a_5396_n6451.n555 6.77231
R5638 a_5396_n6451.n547 a_5396_n6451.t95 5.66511
R5639 a_5396_n6451.n549 a_5396_n6451.n548 5.66379
R5640 a_5396_n6451.n547 a_5396_n6451.n546 5.65285
R5641 a_5396_n6451.n531 a_5396_n6451.n530 5.61877
R5642 a_5396_n6451.n502 a_5396_n6451.t31 5.50607
R5643 a_5396_n6451.n489 a_5396_n6451.t17 5.50607
R5644 a_5396_n6451.n600 a_5396_n6451.t2 5.50607
R5645 a_5396_n6451.n587 a_5396_n6451.t5 5.50607
R5646 a_5396_n6451.n504 a_5396_n6451.n503 5.50475
R5647 a_5396_n6451.n498 a_5396_n6451.n497 5.50475
R5648 a_5396_n6451.n496 a_5396_n6451.t12 5.50475
R5649 a_5396_n6451.n491 a_5396_n6451.n490 5.50475
R5650 a_5396_n6451.n602 a_5396_n6451.n601 5.50475
R5651 a_5396_n6451.n596 a_5396_n6451.n595 5.50475
R5652 a_5396_n6451.n594 a_5396_n6451.t19 5.50475
R5653 a_5396_n6451.n589 a_5396_n6451.n588 5.50475
R5654 a_5396_n6451.n552 a_5396_n6451.n551 4.88835
R5655 a_5396_n6451.n534 a_5396_n6451.n533 4.88517
R5656 a_5396_n6451.n182 a_5396_n6451.n198 1.49912
R5657 a_5396_n6451.n197 a_5396_n6451.n199 1.49876
R5658 a_5396_n6451.n41 a_5396_n6451.n40 1.45673
R5659 a_5396_n6451.n37 a_5396_n6451.n36 1.45673
R5660 a_5396_n6451.n245 a_5396_n6451.n294 2.07625
R5661 a_5396_n6451.n235 a_5396_n6451.n293 2.07625
R5662 a_5396_n6451.n318 a_5396_n6451.n317 2.24588
R5663 a_5396_n6451.n320 a_5396_n6451.n319 2.24588
R5664 a_5396_n6451.n312 a_5396_n6451.n311 2.2453
R5665 a_5396_n6451.n315 a_5396_n6451.n314 2.2453
R5666 a_5396_n6451.n321 a_5396_n6451.n363 4.0312
R5667 a_5396_n6451.n322 a_5396_n6451.n361 5.5012
R5668 a_5396_n6451.n323 a_5396_n6451.t37 5.5012
R5669 a_5396_n6451.n324 a_5396_n6451.n360 4.0312
R5670 a_5396_n6451.n325 a_5396_n6451.n358 5.5012
R5671 a_5396_n6451.n326 a_5396_n6451.t21 5.5012
R5672 a_5396_n6451.n327 a_5396_n6451.n357 4.0312
R5673 a_5396_n6451.n355 a_5396_n6451.n328 5.5012
R5674 a_5396_n6451.t18 a_5396_n6451.n329 5.5012
R5675 a_5396_n6451.n354 a_5396_n6451.n330 4.0312
R5676 a_5396_n6451.n331 a_5396_n6451.n566 4.0312
R5677 a_5396_n6451.n332 a_5396_n6451.n564 5.5012
R5678 a_5396_n6451.n333 a_5396_n6451.t8 5.5012
R5679 a_5396_n6451.n334 a_5396_n6451.n563 4.0312
R5680 a_5396_n6451.n335 a_5396_n6451.n561 5.5012
R5681 a_5396_n6451.n336 a_5396_n6451.t26 5.5012
R5682 a_5396_n6451.n337 a_5396_n6451.n560 4.0312
R5683 a_5396_n6451.n558 a_5396_n6451.n338 5.5012
R5684 a_5396_n6451.t14 a_5396_n6451.n339 5.5012
R5685 a_5396_n6451.n557 a_5396_n6451.n340 4.0312
R5686 a_5396_n6451.n529 a_5396_n6451.n341 4.40099
R5687 a_5396_n6451.n29 a_5396_n6451.n28 0.592804
R5688 a_5396_n6451.n31 a_5396_n6451.n30 0.592804
R5689 a_5396_n6451.n33 a_5396_n6451.n32 0.592804
R5690 a_5396_n6451.n35 a_5396_n6451.n34 0.592804
R5691 a_5396_n6451.n160 a_5396_n6451.n159 0.592738
R5692 a_5396_n6451.n162 a_5396_n6451.n161 0.592738
R5693 a_5396_n6451.n164 a_5396_n6451.n163 0.592738
R5694 a_5396_n6451.n165 a_5396_n6451.n166 0.592738
R5695 a_5396_n6451.n3 a_5396_n6451.n4 0.591918
R5696 a_5396_n6451.n2 a_5396_n6451.n0 0.591918
R5697 a_5396_n6451.n7 a_5396_n6451.n6 0.591918
R5698 a_5396_n6451.n10 a_5396_n6451.n9 0.591918
R5699 a_5396_n6451.n13 a_5396_n6451.n12 0.591918
R5700 a_5396_n6451.n15 a_5396_n6451.n16 0.591918
R5701 a_5396_n6451.n173 a_5396_n6451.n285 1.44185
R5702 a_5396_n6451.n281 a_5396_n6451.n283 1.44185
R5703 a_5396_n6451.n278 a_5396_n6451.n280 1.44185
R5704 a_5396_n6451.n275 a_5396_n6451.n277 1.44185
R5705 a_5396_n6451.n274 a_5396_n6451.n189 1.44185
R5706 a_5396_n6451.n272 a_5396_n6451.n194 1.44185
R5707 a_5396_n6451.n207 a_5396_n6451.n265 1.44113
R5708 a_5396_n6451.n208 a_5396_n6451.n210 1.44113
R5709 a_5396_n6451.n232 a_5396_n6451.n230 1.44113
R5710 a_5396_n6451.n253 a_5396_n6451.n255 1.44113
R5711 a_5396_n6451.n203 a_5396_n6451.n263 1.44113
R5712 a_5396_n6451.n206 a_5396_n6451.n204 1.44113
R5713 a_5396_n6451.n227 a_5396_n6451.n229 1.44113
R5714 a_5396_n6451.n252 a_5396_n6451.n226 1.44113
R5715 a_5396_n6451.n223 a_5396_n6451.n225 1.44113
R5716 a_5396_n6451.n250 a_5396_n6451.n248 1.44113
R5717 a_5396_n6451.n22 a_5396_n6451.n21 0.604258
R5718 a_5396_n6451.n211 a_5396_n6451.n233 1.44113
R5719 a_5396_n6451.n6 a_5396_n6451.n8 0.591264
R5720 a_5396_n6451.n177 a_5396_n6451.n178 1.44113
R5721 a_5396_n6451.n282 a_5396_n6451.n281 1.44113
R5722 a_5396_n6451.n0 a_5396_n6451.n1 0.591264
R5723 a_5396_n6451.n174 a_5396_n6451.n176 1.44113
R5724 a_5396_n6451.n173 a_5396_n6451.n284 1.44113
R5725 a_5396_n6451.n5 a_5396_n6451.n3 0.591264
R5726 a_5396_n6451.n172 a_5396_n6451.n171 0.0478472
R5727 a_5396_n6451.n181 a_5396_n6451.n182 1.44113
R5728 a_5396_n6451.n279 a_5396_n6451.n278 1.44113
R5729 a_5396_n6451.n198 a_5396_n6451.n180 0.0193886
R5730 a_5396_n6451.n183 a_5396_n6451.n181 1.44113
R5731 a_5396_n6451.n179 a_5396_n6451.n177 1.44113
R5732 a_5396_n6451.n174 a_5396_n6451.n175 1.44113
R5733 a_5396_n6451.n269 a_5396_n6451.n218 1.44113
R5734 a_5396_n6451.n221 a_5396_n6451.n219 1.44113
R5735 a_5396_n6451.n244 a_5396_n6451.n217 1.44113
R5736 a_5396_n6451.n242 a_5396_n6451.n262 1.44113
R5737 a_5396_n6451.n267 a_5396_n6451.n213 1.44113
R5738 a_5396_n6451.n216 a_5396_n6451.n214 1.44113
R5739 a_5396_n6451.n241 a_5396_n6451.n212 1.44113
R5740 a_5396_n6451.n239 a_5396_n6451.n260 1.44113
R5741 a_5396_n6451.n238 a_5396_n6451.n236 1.44113
R5742 a_5396_n6451.n256 a_5396_n6451.n258 1.44113
R5743 a_5396_n6451.n19 a_5396_n6451.n18 0.604258
R5744 a_5396_n6451.n222 a_5396_n6451.n247 1.44113
R5745 a_5396_n6451.n294 a_5396_n6451.n246 0.0221358
R5746 a_5396_n6451.n222 a_5396_n6451.n245 1.44113
R5747 a_5396_n6451.n18 a_5396_n6451.n20 0.604258
R5748 a_5396_n6451.n261 a_5396_n6451.n242 1.44113
R5749 a_5396_n6451.n217 a_5396_n6451.n243 1.44113
R5750 a_5396_n6451.n219 a_5396_n6451.n220 1.44113
R5751 a_5396_n6451.n218 a_5396_n6451.n270 1.44113
R5752 a_5396_n6451.n259 a_5396_n6451.n239 1.44113
R5753 a_5396_n6451.n212 a_5396_n6451.n240 1.44113
R5754 a_5396_n6451.n214 a_5396_n6451.n215 1.44113
R5755 a_5396_n6451.n213 a_5396_n6451.n268 1.44113
R5756 a_5396_n6451.n257 a_5396_n6451.n256 1.44113
R5757 a_5396_n6451.n237 a_5396_n6451.n236 1.44113
R5758 a_5396_n6451.n24 a_5396_n6451.n25 0.0301596
R5759 a_5396_n6451.n17 a_5396_n6451.n15 0.591264
R5760 a_5396_n6451.n192 a_5396_n6451.n190 1.44113
R5761 a_5396_n6451.n189 a_5396_n6451.n273 1.44113
R5762 a_5396_n6451.n12 a_5396_n6451.n14 0.591264
R5763 a_5396_n6451.n186 a_5396_n6451.n187 1.44113
R5764 a_5396_n6451.n276 a_5396_n6451.n275 1.44113
R5765 a_5396_n6451.n9 a_5396_n6451.n11 0.591264
R5766 a_5396_n6451.n184 a_5396_n6451.n185 0.0478472
R5767 a_5396_n6451.n197 a_5396_n6451.n195 1.44113
R5768 a_5396_n6451.n194 a_5396_n6451.n271 1.44113
R5769 a_5396_n6451.n193 a_5396_n6451.n199 0.0193886
R5770 a_5396_n6451.n195 a_5396_n6451.n196 1.44113
R5771 a_5396_n6451.n190 a_5396_n6451.n191 1.44113
R5772 a_5396_n6451.n188 a_5396_n6451.n186 1.44113
R5773 a_5396_n6451.n234 a_5396_n6451.n293 0.0221358
R5774 a_5396_n6451.n235 a_5396_n6451.n211 1.44113
R5775 a_5396_n6451.n21 a_5396_n6451.n23 0.604258
R5776 a_5396_n6451.n254 a_5396_n6451.n253 1.44113
R5777 a_5396_n6451.n231 a_5396_n6451.n230 1.44113
R5778 a_5396_n6451.n208 a_5396_n6451.n209 1.44113
R5779 a_5396_n6451.n266 a_5396_n6451.n207 1.44113
R5780 a_5396_n6451.n226 a_5396_n6451.n251 1.44113
R5781 a_5396_n6451.n228 a_5396_n6451.n227 1.44113
R5782 a_5396_n6451.n205 a_5396_n6451.n204 1.44113
R5783 a_5396_n6451.n264 a_5396_n6451.n203 1.44113
R5784 a_5396_n6451.n248 a_5396_n6451.n249 1.44113
R5785 a_5396_n6451.n223 a_5396_n6451.n224 1.44113
R5786 a_5396_n6451.n26 a_5396_n6451.n27 0.0301596
R5787 a_5396_n6451.n392 a_5396_n6451.n391 4.5005
R5788 a_5396_n6451.n153 a_5396_n6451.n152 2.21666
R5789 a_5396_n6451.n394 a_5396_n6451.n393 4.5005
R5790 a_5396_n6451.n108 a_5396_n6451.n390 4.5005
R5791 a_5396_n6451.n109 a_5396_n6451.n110 2.21666
R5792 a_5396_n6451.n123 a_5396_n6451.n122 2.21666
R5793 a_5396_n6451.n398 a_5396_n6451.n389 4.5005
R5794 a_5396_n6451.n137 a_5396_n6451.n136 2.21666
R5795 a_5396_n6451.n400 a_5396_n6451.n399 4.5005
R5796 a_5396_n6451.n156 a_5396_n6451.n154 2.21666
R5797 a_5396_n6451.n401 a_5396_n6451.n155 4.5005
R5798 a_5396_n6451.n316 a_5396_n6451.n402 4.5005
R5799 a_5396_n6451.n404 a_5396_n6451.n403 4.5005
R5800 a_5396_n6451.n140 a_5396_n6451.n138 2.21666
R5801 a_5396_n6451.n405 a_5396_n6451.n139 4.5005
R5802 a_5396_n6451.n157 a_5396_n6451.n158 2.21666
R5803 a_5396_n6451.n407 a_5396_n6451.n406 4.5005
R5804 a_5396_n6451.n112 a_5396_n6451.n114 4.5005
R5805 a_5396_n6451.n115 a_5396_n6451.n113 2.21666
R5806 a_5396_n6451.n126 a_5396_n6451.n125 2.21666
R5807 a_5396_n6451.n124 a_5396_n6451.n412 4.5005
R5808 a_5396_n6451.n143 a_5396_n6451.n142 2.21666
R5809 a_5396_n6451.n141 a_5396_n6451.n411 4.5005
R5810 a_5396_n6451.n167 a_5396_n6451.n168 0.332154
R5811 a_5396_n6451.n48 a_5396_n6451.n46 2.21666
R5812 a_5396_n6451.n45 a_5396_n6451.n47 4.5005
R5813 a_5396_n6451.n51 a_5396_n6451.n50 2.21666
R5814 a_5396_n6451.n49 a_5396_n6451.n382 4.5005
R5815 a_5396_n6451.n381 a_5396_n6451.n378 4.5005
R5816 a_5396_n6451.n432 a_5396_n6451.n431 4.5005
R5817 a_5396_n6451.n58 a_5396_n6451.n59 2.21666
R5818 a_5396_n6451.n430 a_5396_n6451.n56 4.5005
R5819 a_5396_n6451.n57 a_5396_n6451.n55 2.21666
R5820 a_5396_n6451.n429 a_5396_n6451.n54 4.5005
R5821 a_5396_n6451.n53 a_5396_n6451.n52 2.21666
R5822 a_5396_n6451.n61 a_5396_n6451.n60 2.21666
R5823 a_5396_n6451.n422 a_5396_n6451.n388 4.5005
R5824 a_5396_n6451.n63 a_5396_n6451.n62 2.21666
R5825 a_5396_n6451.n423 a_5396_n6451.n387 4.5005
R5826 a_5396_n6451.n65 a_5396_n6451.n64 2.21666
R5827 a_5396_n6451.n425 a_5396_n6451.n424 4.5005
R5828 a_5396_n6451.n426 a_5396_n6451.n386 4.5005
R5829 a_5396_n6451.n418 a_5396_n6451.n417 4.5005
R5830 a_5396_n6451.n69 a_5396_n6451.n68 2.21666
R5831 a_5396_n6451.n416 a_5396_n6451.n415 4.5005
R5832 a_5396_n6451.n67 a_5396_n6451.n66 2.21666
R5833 a_5396_n6451.n39 a_5396_n6451.n38 0.349872
R5834 a_5396_n6451.n434 a_5396_n6451.n309 4.5005
R5835 a_5396_n6451.n144 a_5396_n6451.n145 2.21666
R5836 a_5396_n6451.n436 a_5396_n6451.n435 4.5005
R5837 a_5396_n6451.n102 a_5396_n6451.n104 4.5005
R5838 a_5396_n6451.n105 a_5396_n6451.n103 2.21666
R5839 a_5396_n6451.n118 a_5396_n6451.n117 2.21666
R5840 a_5396_n6451.n116 a_5396_n6451.n455 4.5005
R5841 a_5396_n6451.n129 a_5396_n6451.n128 2.21666
R5842 a_5396_n6451.n127 a_5396_n6451.n440 4.5005
R5843 a_5396_n6451.n147 a_5396_n6451.n148 2.21666
R5844 a_5396_n6451.n146 a_5396_n6451.n441 4.5005
R5845 a_5396_n6451.n454 a_5396_n6451.n453 4.5005
R5846 a_5396_n6451.n313 a_5396_n6451.n452 4.5005
R5847 a_5396_n6451.n132 a_5396_n6451.n131 2.21666
R5848 a_5396_n6451.n130 a_5396_n6451.n442 4.5005
R5849 a_5396_n6451.n150 a_5396_n6451.n151 2.21666
R5850 a_5396_n6451.n149 a_5396_n6451.n443 4.5005
R5851 a_5396_n6451.n451 a_5396_n6451.n450 4.5005
R5852 a_5396_n6451.n107 a_5396_n6451.n106 2.21666
R5853 a_5396_n6451.n120 a_5396_n6451.n121 2.21666
R5854 a_5396_n6451.n119 a_5396_n6451.n445 4.5005
R5855 a_5396_n6451.n134 a_5396_n6451.n135 2.21666
R5856 a_5396_n6451.n133 a_5396_n6451.n446 4.5005
R5857 a_5396_n6451.n169 a_5396_n6451.n170 0.332154
R5858 a_5396_n6451.n71 a_5396_n6451.n72 2.21666
R5859 a_5396_n6451.n70 a_5396_n6451.n371 4.5005
R5860 a_5396_n6451.n74 a_5396_n6451.n75 2.21666
R5861 a_5396_n6451.n73 a_5396_n6451.n372 4.5005
R5862 a_5396_n6451.n376 a_5396_n6451.n375 4.5005
R5863 a_5396_n6451.n82 a_5396_n6451.n370 4.5005
R5864 a_5396_n6451.n83 a_5396_n6451.n84 2.21666
R5865 a_5396_n6451.n79 a_5396_n6451.n369 4.5005
R5866 a_5396_n6451.n80 a_5396_n6451.n81 2.21666
R5867 a_5396_n6451.n76 a_5396_n6451.n368 4.5005
R5868 a_5396_n6451.n78 a_5396_n6451.n77 2.21666
R5869 a_5396_n6451.n89 a_5396_n6451.n87 2.21666
R5870 a_5396_n6451.n86 a_5396_n6451.n88 4.5005
R5871 a_5396_n6451.n92 a_5396_n6451.n91 2.21666
R5872 a_5396_n6451.n90 a_5396_n6451.n476 4.5005
R5873 a_5396_n6451.n95 a_5396_n6451.n94 2.21666
R5874 a_5396_n6451.n93 a_5396_n6451.n366 4.5005
R5875 a_5396_n6451.n475 a_5396_n6451.n474 4.5005
R5876 a_5396_n6451.n482 a_5396_n6451.n481 4.5005
R5877 a_5396_n6451.n99 a_5396_n6451.n100 2.21666
R5878 a_5396_n6451.n480 a_5396_n6451.n97 4.5005
R5879 a_5396_n6451.n98 a_5396_n6451.n96 2.21666
R5880 a_5396_n6451.n42 a_5396_n6451.n43 0.349872
R5881 a_5396_n6451.n537 a_5396_n6451.n536 4.40142
R5882 a_5396_n6451.n348 a_5396_n6451.n347 4.24002
R5883 a_5396_n6451.n345 a_5396_n6451.n344 4.24002
R5884 a_5396_n6451.n574 a_5396_n6451.n573 4.24002
R5885 a_5396_n6451.n520 a_5396_n6451.n519 4.24002
R5886 a_5396_n6451.n507 a_5396_n6451.n506 4.03475
R5887 a_5396_n6451.n501 a_5396_n6451.n500 4.03475
R5888 a_5396_n6451.n495 a_5396_n6451.n494 4.03475
R5889 a_5396_n6451.n488 a_5396_n6451.n487 4.03475
R5890 a_5396_n6451.n605 a_5396_n6451.n604 4.03475
R5891 a_5396_n6451.n599 a_5396_n6451.n598 4.03475
R5892 a_5396_n6451.n593 a_5396_n6451.n592 4.03475
R5893 a_5396_n6451.n586 a_5396_n6451.n585 4.03475
R5894 a_5396_n6451.n537 a_5396_n6451.n535 3.84721
R5895 a_5396_n6451.n348 a_5396_n6451.n346 3.68818
R5896 a_5396_n6451.n345 a_5396_n6451.n343 3.68818
R5897 a_5396_n6451.n574 a_5396_n6451.n572 3.68818
R5898 a_5396_n6451.n520 a_5396_n6451.n518 3.68818
R5899 a_5396_n6451.n554 a_5396_n6451.n517 3.48654
R5900 a_5396_n6451.n569 a_5396_n6451.n554 3.42822
R5901 a_5396_n6451.n466 a_5396_n6451.n364 3.37173
R5902 a_5396_n6451.n582 a_5396_n6451.n581 3.23904
R5903 a_5396_n6451.n516 a_5396_n6451.n515 3.23904
R5904 a_5396_n6451.n544 a_5396_n6451.n543 3.23004
R5905 a_5396_n6451.n542 a_5396_n6451.n541 3.14142
R5906 a_5396_n6451.n514 a_5396_n6451.n513 2.77002
R5907 a_5396_n6451.n580 a_5396_n6451.n579 2.77002
R5908 a_5396_n6451.n525 a_5396_n6451.n524 2.77002
R5909 a_5396_n6451.n618 a_5396_n6451.n617 2.77002
R5910 a_5396_n6451.n614 a_5396_n6451.n345 2.7375
R5911 a_5396_n6451.n526 a_5396_n6451.n520 2.73714
R5912 a_5396_n6451.n543 a_5396_n6451.n537 2.71914
R5913 a_5396_n6451.n498 a_5396_n6451.n496 2.60203
R5914 a_5396_n6451.n596 a_5396_n6451.n594 2.60203
R5915 a_5396_n6451.n542 a_5396_n6451.n539 2.58721
R5916 a_5396_n6451.n549 a_5396_n6451.n547 2.55136
R5917 a_5396_n6451.n491 a_5396_n6451.n489 2.52436
R5918 a_5396_n6451.n504 a_5396_n6451.n502 2.52436
R5919 a_5396_n6451.n589 a_5396_n6451.n587 2.52436
R5920 a_5396_n6451.n602 a_5396_n6451.n600 2.52436
R5921 a_5396_n6451.n198 a_5396_n6451.n183 1.48408
R5922 a_5396_n6451.n196 a_5396_n6451.n199 1.48372
R5923 a_5396_n6451.n467 a_5396_n6451.n465 2.40699
R5924 a_5396_n6451.n433 a_5396_n6451.n377 2.30989
R5925 a_5396_n6451.n413 a_5396_n6451.n111 2.30989
R5926 a_5396_n6451.n544 a_5396_n6451.n534 2.2807
R5927 a_5396_n6451.n473 a_5396_n6451.n367 2.25752
R5928 a_5396_n6451.n428 a_5396_n6451.n427 2.25752
R5929 a_5396_n6451.n289 a_5396_n6451.n288 1.44642
R5930 a_5396_n6451.n290 a_5396_n6451.n200 1.44642
R5931 a_5396_n6451.n291 a_5396_n6451.n201 1.44642
R5932 a_5396_n6451.n292 a_5396_n6451.n202 1.44642
R5933 a_5396_n6451.n301 a_5396_n6451.n300 1.44612
R5934 a_5396_n6451.n302 a_5396_n6451.n286 1.44612
R5935 a_5396_n6451.n303 a_5396_n6451.n287 1.44612
R5936 a_5396_n6451.n305 a_5396_n6451.n304 1.44612
R5937 a_5396_n6451.n514 a_5396_n6451.n511 2.21818
R5938 a_5396_n6451.n580 a_5396_n6451.n577 2.21818
R5939 a_5396_n6451.n525 a_5396_n6451.n522 2.21818
R5940 a_5396_n6451.n617 a_5396_n6451.n616 2.21818
R5941 a_5396_n6451.n261 a_5396_n6451.n459 2.23847
R5942 a_5396_n6451.n298 a_5396_n6451.n257 2.23847
R5943 a_5396_n6451.n299 a_5396_n6451.n254 2.23847
R5944 a_5396_n6451.n249 a_5396_n6451.n464 2.23847
R5945 a_5396_n6451.n458 a_5396_n6451.n296 2.07182
R5946 a_5396_n6451.n460 a_5396_n6451.n295 2.07182
R5947 a_5396_n6451.n296 a_5396_n6451.n7 2.46476
R5948 a_5396_n6451.n4 a_5396_n6451.n295 2.46476
R5949 a_5396_n6451.n16 a_5396_n6451.n461 2.46476
R5950 a_5396_n6451.n297 a_5396_n6451.n10 2.46476
R5951 a_5396_n6451.n463 a_5396_n6451.n364 1.80314
R5952 a_5396_n6451.n571 a_5396_n6451.n526 1.73904
R5953 a_5396_n6451.n614 a_5396_n6451.n613 1.73868
R5954 a_5396_n6451.n509 a_5396_n6451.n484 1.70908
R5955 a_5396_n6451.n468 a_5396_n6451.n467 1.68395
R5956 a_5396_n6451.n484 a_5396_n6451.n483 1.68395
R5957 a_5396_n6451.n461 a_5396_n6451.n457 1.5005
R5958 a_5396_n6451.n459 a_5396_n6451.n458 1.5005
R5959 a_5396_n6451.n465 a_5396_n6451.n299 1.5005
R5960 a_5396_n6451.n464 a_5396_n6451.n463 1.5005
R5961 a_5396_n6451.n462 a_5396_n6451.n297 1.5005
R5962 a_5396_n6451.n460 a_5396_n6451.n298 1.5005
R5963 a_5396_n6451.n456 a_5396_n6451.n101 1.5005
R5964 a_5396_n6451.n433 a_5396_n6451.n44 1.5005
R5965 a_5396_n6451.n469 a_5396_n6451.n468 1.5005
R5966 a_5396_n6451.n483 a_5396_n6451.n85 1.5005
R5967 a_5396_n6451.n444 a_5396_n6451.n365 1.5005
R5968 a_5396_n6451.n414 a_5396_n6451.n413 1.5005
R5969 a_5396_n6451.n569 a_5396_n6451.n568 1.5005
R5970 a_5396_n6451.n571 a_5396_n6451.n570 1.5005
R5971 a_5396_n6451.n590 a_5396_n6451.n351 1.5005
R5972 a_5396_n6451.n611 a_5396_n6451.n610 1.5005
R5973 a_5396_n6451.n492 a_5396_n6451.n350 1.5005
R5974 a_5396_n6451.n553 a_5396_n6451.n552 1.5005
R5975 a_5396_n6451.n567 a_5396_n6451.n517 1.5005
R5976 a_5396_n6451.n607 a_5396_n6451.n606 1.5005
R5977 a_5396_n6451.n609 a_5396_n6451.n608 1.5005
R5978 a_5396_n6451.n509 a_5396_n6451.n508 1.5005
R5979 a_5396_n6451.n613 a_5396_n6451.n612 1.5005
R5980 a_5396_n6451.n458 a_5396_n6451.n457 1.47516
R5981 a_5396_n6451.n462 a_5396_n6451.n460 1.47516
R5982 a_5396_n6451.n616 a_5396_n6451.t40 1.4705
R5983 a_5396_n6451.n616 a_5396_n6451.n615 1.4705
R5984 a_5396_n6451.n511 a_5396_n6451.t22 1.4705
R5985 a_5396_n6451.n511 a_5396_n6451.n510 1.4705
R5986 a_5396_n6451.n513 a_5396_n6451.t23 1.4705
R5987 a_5396_n6451.n513 a_5396_n6451.n512 1.4705
R5988 a_5396_n6451.n506 a_5396_n6451.t11 1.4705
R5989 a_5396_n6451.n506 a_5396_n6451.n505 1.4705
R5990 a_5396_n6451.n500 a_5396_n6451.t24 1.4705
R5991 a_5396_n6451.n500 a_5396_n6451.n499 1.4705
R5992 a_5396_n6451.n494 a_5396_n6451.t3 1.4705
R5993 a_5396_n6451.n494 a_5396_n6451.n493 1.4705
R5994 a_5396_n6451.n487 a_5396_n6451.t38 1.4705
R5995 a_5396_n6451.n487 a_5396_n6451.n486 1.4705
R5996 a_5396_n6451.n363 a_5396_n6451.t10 1.4705
R5997 a_5396_n6451.n363 a_5396_n6451.n362 1.4705
R5998 a_5396_n6451.n360 a_5396_n6451.t7 1.4705
R5999 a_5396_n6451.n360 a_5396_n6451.n359 1.4705
R6000 a_5396_n6451.n357 a_5396_n6451.t28 1.4705
R6001 a_5396_n6451.n357 a_5396_n6451.n356 1.4705
R6002 a_5396_n6451.n354 a_5396_n6451.t15 1.4705
R6003 a_5396_n6451.n354 a_5396_n6451.n353 1.4705
R6004 a_5396_n6451.n604 a_5396_n6451.t6 1.4705
R6005 a_5396_n6451.n604 a_5396_n6451.n603 1.4705
R6006 a_5396_n6451.n598 a_5396_n6451.t27 1.4705
R6007 a_5396_n6451.n598 a_5396_n6451.n597 1.4705
R6008 a_5396_n6451.n592 a_5396_n6451.t4 1.4705
R6009 a_5396_n6451.n592 a_5396_n6451.n591 1.4705
R6010 a_5396_n6451.n585 a_5396_n6451.t25 1.4705
R6011 a_5396_n6451.n585 a_5396_n6451.n584 1.4705
R6012 a_5396_n6451.n577 a_5396_n6451.t33 1.4705
R6013 a_5396_n6451.n577 a_5396_n6451.n576 1.4705
R6014 a_5396_n6451.n579 a_5396_n6451.t32 1.4705
R6015 a_5396_n6451.n579 a_5396_n6451.n578 1.4705
R6016 a_5396_n6451.n522 a_5396_n6451.t36 1.4705
R6017 a_5396_n6451.n522 a_5396_n6451.n521 1.4705
R6018 a_5396_n6451.n524 a_5396_n6451.t35 1.4705
R6019 a_5396_n6451.n524 a_5396_n6451.n523 1.4705
R6020 a_5396_n6451.n566 a_5396_n6451.t16 1.4705
R6021 a_5396_n6451.n566 a_5396_n6451.n565 1.4705
R6022 a_5396_n6451.n563 a_5396_n6451.t34 1.4705
R6023 a_5396_n6451.n563 a_5396_n6451.n562 1.4705
R6024 a_5396_n6451.n560 a_5396_n6451.t9 1.4705
R6025 a_5396_n6451.n560 a_5396_n6451.n559 1.4705
R6026 a_5396_n6451.n557 a_5396_n6451.t29 1.4705
R6027 a_5396_n6451.n557 a_5396_n6451.n556 1.4705
R6028 a_5396_n6451.t41 a_5396_n6451.n618 1.4705
R6029 a_5396_n6451.n618 a_5396_n6451.n342 1.4705
R6030 a_5396_n6451.n515 a_5396_n6451.n514 1.46537
R6031 a_5396_n6451.n349 a_5396_n6451.n348 1.46537
R6032 a_5396_n6451.n581 a_5396_n6451.n580 1.46537
R6033 a_5396_n6451.n575 a_5396_n6451.n574 1.46537
R6034 a_5396_n6451.n526 a_5396_n6451.n525 1.46537
R6035 a_5396_n6451.n543 a_5396_n6451.n542 1.46537
R6036 a_5396_n6451.n617 a_5396_n6451.n614 1.46537
R6037 a_5396_n6451.n554 a_5396_n6451.n553 1.41182
R6038 a_5396_n6451.n307 a_5396_n6451.t281 8.40801
R6039 a_5396_n6451.n308 a_5396_n6451.t206 8.40801
R6040 a_5396_n6451.n496 a_5396_n6451.n495 1.27228
R6041 a_5396_n6451.n501 a_5396_n6451.n498 1.27228
R6042 a_5396_n6451.n594 a_5396_n6451.n593 1.27228
R6043 a_5396_n6451.n599 a_5396_n6451.n596 1.27228
R6044 a_5396_n6451.n581 a_5396_n6451.n575 1.27228
R6045 a_5396_n6451.n515 a_5396_n6451.n349 1.27228
R6046 a_5396_n6451.n489 a_5396_n6451.n488 1.26756
R6047 a_5396_n6451.n502 a_5396_n6451.n501 1.26756
R6048 a_5396_n6451.n587 a_5396_n6451.n586 1.26756
R6049 a_5396_n6451.n600 a_5396_n6451.n599 1.26756
R6050 a_5396_n6451.n551 a_5396_n6451.t0 1.2605
R6051 a_5396_n6451.n551 a_5396_n6451.n550 1.2605
R6052 a_5396_n6451.n546 a_5396_n6451.t1 1.2605
R6053 a_5396_n6451.n546 a_5396_n6451.n545 1.2605
R6054 a_5396_n6451.n539 a_5396_n6451.t91 1.2605
R6055 a_5396_n6451.n539 a_5396_n6451.n538 1.2605
R6056 a_5396_n6451.n541 a_5396_n6451.t104 1.2605
R6057 a_5396_n6451.n541 a_5396_n6451.n540 1.2605
R6058 a_5396_n6451.n533 a_5396_n6451.t99 1.2605
R6059 a_5396_n6451.n533 a_5396_n6451.n532 1.2605
R6060 a_5396_n6451.n529 a_5396_n6451.t96 1.2605
R6061 a_5396_n6451.n529 a_5396_n6451.n528 1.2605
R6062 a_5396_n6451.n125 a_5396_n6451.n410 1.24866
R6063 a_5396_n6451.n122 a_5396_n6451.n397 1.24866
R6064 a_5396_n6451.n447 a_5396_n6451.n120 1.24866
R6065 a_5396_n6451.n117 a_5396_n6451.n439 1.24866
R6066 a_5396_n6451.n408 a_5396_n6451.n115 1.24629
R6067 a_5396_n6451.n395 a_5396_n6451.n109 1.24629
R6068 a_5396_n6451.n106 a_5396_n6451.n449 1.24629
R6069 a_5396_n6451.n437 a_5396_n6451.n105 1.24629
R6070 a_5396_n6451.n456 a_5396_n6451.n433 1.23709
R6071 a_5396_n6451.n413 a_5396_n6451.n365 1.23709
R6072 a_5396_n6451.n477 a_5396_n6451.n89 1.22261
R6073 a_5396_n6451.n470 a_5396_n6451.n71 1.22261
R6074 a_5396_n6451.n60 a_5396_n6451.n421 1.22261
R6075 a_5396_n6451.n383 a_5396_n6451.n48 1.22261
R6076 a_5396_n6451.n481 a_5396_n6451.n479 1.21313
R6077 a_5396_n6451.n82 a_5396_n6451.n472 1.21313
R6078 a_5396_n6451.n419 a_5396_n6451.n418 1.21313
R6079 a_5396_n6451.n431 a_5396_n6451.n385 1.21313
R6080 a_5396_n6451.n381 a_5396_n6451.n380 1.12904
R6081 a_5396_n6451.n375 a_5396_n6451.n374 1.12904
R6082 a_5396_n6451.n466 a_5396_n6451.n350 1.10472
R6083 a_5396_n6451.n468 a_5396_n6451.n456 0.809892
R6084 a_5396_n6451.n483 a_5396_n6451.n365 0.809892
R6085 a_5396_n6451.n492 a_5396_n6451.n491 0.796291
R6086 a_5396_n6451.n508 a_5396_n6451.n504 0.796291
R6087 a_5396_n6451.n590 a_5396_n6451.n589 0.796291
R6088 a_5396_n6451.n606 a_5396_n6451.n602 0.796291
R6089 a_5396_n6451.n612 a_5396_n6451.n611 0.780703
R6090 a_5396_n6451.n570 a_5396_n6451.n569 0.780703
R6091 a_5396_n6451.n608 a_5396_n6451.n516 0.780703
R6092 a_5396_n6451.n582 a_5396_n6451.n517 0.780703
R6093 a_5396_n6451.n552 a_5396_n6451.n549 0.769291
R6094 a_5396_n6451.n534 a_5396_n6451.n531 0.767125
R6095 a_5396_n6451.n123 a_5396_n6451.n377 0.821185
R6096 a_5396_n6451.n111 a_5396_n6451.n126 0.821185
R6097 a_5396_n6451.n101 a_5396_n6451.n118 0.821185
R6098 a_5396_n6451.n121 a_5396_n6451.n444 0.821185
R6099 a_5396_n6451.n44 a_5396_n6451.n432 0.71825
R6100 a_5396_n6451.n417 a_5396_n6451.n414 0.71825
R6101 a_5396_n6451.n469 a_5396_n6451.n370 0.71825
R6102 a_5396_n6451.n85 a_5396_n6451.n482 0.71825
R6103 a_5396_n6451.n478 a_5396_n6451.n477 0.673132
R6104 a_5396_n6451.n479 a_5396_n6451.n478 0.673132
R6105 a_5396_n6451.n471 a_5396_n6451.n470 0.673132
R6106 a_5396_n6451.n472 a_5396_n6451.n471 0.673132
R6107 a_5396_n6451.n409 a_5396_n6451.n408 0.673132
R6108 a_5396_n6451.n410 a_5396_n6451.n409 0.673132
R6109 a_5396_n6451.n396 a_5396_n6451.n395 0.673132
R6110 a_5396_n6451.n397 a_5396_n6451.n396 0.673132
R6111 a_5396_n6451.n421 a_5396_n6451.n420 0.673132
R6112 a_5396_n6451.n420 a_5396_n6451.n419 0.673132
R6113 a_5396_n6451.n384 a_5396_n6451.n383 0.673132
R6114 a_5396_n6451.n385 a_5396_n6451.n384 0.673132
R6115 a_5396_n6451.n449 a_5396_n6451.n448 0.673132
R6116 a_5396_n6451.n448 a_5396_n6451.n447 0.673132
R6117 a_5396_n6451.n438 a_5396_n6451.n437 0.673132
R6118 a_5396_n6451.n439 a_5396_n6451.n438 0.673132
R6119 a_5396_n6451.n612 a_5396_n6451.n350 0.638405
R6120 a_5396_n6451.n570 a_5396_n6451.n351 0.638405
R6121 a_5396_n6451.n553 a_5396_n6451.n544 0.638405
R6122 a_5396_n6451.n516 a_5396_n6451.n509 0.638405
R6123 a_5396_n6451.n607 a_5396_n6451.n582 0.638405
R6124 a_5396_n6451.n611 a_5396_n6451.n351 0.628372
R6125 a_5396_n6451.n608 a_5396_n6451.n607 0.628372
R6126 a_5396_n6451.n484 a_5396_n6451.n364 0.604355
R6127 a_5396_n6451.n467 a_5396_n6451.n466 0.603852
R6128 a_5396_n6451.n465 a_5396_n6451.n457 0.571818
R6129 a_5396_n6451.n463 a_5396_n6451.n462 0.571818
R6130 a_5396_n6451.n495 a_5396_n6451.n492 0.476484
R6131 a_5396_n6451.n508 a_5396_n6451.n507 0.476484
R6132 a_5396_n6451.n593 a_5396_n6451.n590 0.476484
R6133 a_5396_n6451.n606 a_5396_n6451.n605 0.476484
R6134 a_5396_n6451.n307 a_5396_n6451.n306 0.307602
R6135 a_5396_n6451.n310 a_5396_n6451.n308 0.307602
R6136 a_5396_n6451.n141 a_5396_n6451.n167 0.394842
R6137 a_5396_n6451.n157 a_5396_n6451.n139 0.394842
R6138 a_5396_n6451.n156 a_5396_n6451.n400 0.394842
R6139 a_5396_n6451.n152 a_5396_n6451.n392 0.394842
R6140 a_5396_n6451.n133 a_5396_n6451.n169 0.394842
R6141 a_5396_n6451.n130 a_5396_n6451.n150 0.394842
R6142 a_5396_n6451.n127 a_5396_n6451.n147 0.394842
R6143 a_5396_n6451.n144 a_5396_n6451.n309 0.394842
R6144 a_5396_n6451.n124 a_5396_n6451.n142 0.381816
R6145 a_5396_n6451.n140 a_5396_n6451.n404 0.381816
R6146 a_5396_n6451.n136 a_5396_n6451.n398 0.381816
R6147 a_5396_n6451.n119 a_5396_n6451.n134 0.381816
R6148 a_5396_n6451.n313 a_5396_n6451.n131 0.381816
R6149 a_5396_n6451.n116 a_5396_n6451.n128 0.381816
R6150 a_5396_n6451.n99 a_5396_n6451.n97 0.379447
R6151 a_5396_n6451.n98 a_5396_n6451.n42 0.379447
R6152 a_5396_n6451.n93 a_5396_n6451.n475 0.379447
R6153 a_5396_n6451.n90 a_5396_n6451.n94 0.379447
R6154 a_5396_n6451.n91 a_5396_n6451.n88 0.379447
R6155 a_5396_n6451.n79 a_5396_n6451.n83 0.379447
R6156 a_5396_n6451.n76 a_5396_n6451.n80 0.379447
R6157 a_5396_n6451.n73 a_5396_n6451.n376 0.379447
R6158 a_5396_n6451.n70 a_5396_n6451.n74 0.379447
R6159 a_5396_n6451.n68 a_5396_n6451.n416 0.379447
R6160 a_5396_n6451.n66 a_5396_n6451.n39 0.379447
R6161 a_5396_n6451.n426 a_5396_n6451.n425 0.379447
R6162 a_5396_n6451.n64 a_5396_n6451.n423 0.379447
R6163 a_5396_n6451.n62 a_5396_n6451.n422 0.379447
R6164 a_5396_n6451.n58 a_5396_n6451.n56 0.379447
R6165 a_5396_n6451.n57 a_5396_n6451.n429 0.379447
R6166 a_5396_n6451.n49 a_5396_n6451.n378 0.379447
R6167 a_5396_n6451.n50 a_5396_n6451.n47 0.379447
R6168 a_5396_n6451.n210 a_5396_n6451.n232 0.647707
R6169 a_5396_n6451.n206 a_5396_n6451.n229 0.647707
R6170 a_5396_n6451.n27 a_5396_n6451.n225 1.48545
R6171 a_5396_n6451.n178 a_5396_n6451.n8 0.908313
R6172 a_5396_n6451.n5 a_5396_n6451.n172 1.74614
R6173 a_5396_n6451.n221 a_5396_n6451.n244 0.647707
R6174 a_5396_n6451.n216 a_5396_n6451.n241 0.647707
R6175 a_5396_n6451.n25 a_5396_n6451.n238 1.48545
R6176 a_5396_n6451.n220 a_5396_n6451.n243 0.647707
R6177 a_5396_n6451.n215 a_5396_n6451.n240 0.647707
R6178 a_5396_n6451.n25 a_5396_n6451.n237 1.48641
R6179 a_5396_n6451.n192 a_5396_n6451.n17 0.907953
R6180 a_5396_n6451.n14 a_5396_n6451.n187 0.908313
R6181 a_5396_n6451.n185 a_5396_n6451.n11 1.74614
R6182 a_5396_n6451.n209 a_5396_n6451.n231 0.647707
R6183 a_5396_n6451.n228 a_5396_n6451.n205 0.647707
R6184 a_5396_n6451.n27 a_5396_n6451.n224 1.48641
R6185 a_5396_n6451.n153 a_5396_n6451.n391 0.44431
R6186 a_5396_n6451.n399 a_5396_n6451.n154 0.44431
R6187 a_5396_n6451.n158 a_5396_n6451.n405 0.44431
R6188 a_5396_n6451.n168 a_5396_n6451.n411 1.20531
R6189 a_5396_n6451.n145 a_5396_n6451.n434 0.44431
R6190 a_5396_n6451.n148 a_5396_n6451.n440 0.44431
R6191 a_5396_n6451.n151 a_5396_n6451.n442 0.44431
R6192 a_5396_n6451.n170 a_5396_n6451.n446 1.20531
R6193 a_5396_n6451.n233 a_5396_n6451.n293 2.07535
R6194 a_5396_n6451.n232 a_5396_n6451.n255 0.635332
R6195 a_5396_n6451.n229 a_5396_n6451.n252 0.635332
R6196 a_5396_n6451.n225 a_5396_n6451.n250 0.635332
R6197 a_5396_n6451.n247 a_5396_n6451.n294 2.07535
R6198 a_5396_n6451.n244 a_5396_n6451.n262 0.635332
R6199 a_5396_n6451.n241 a_5396_n6451.n260 0.635332
R6200 a_5396_n6451.n238 a_5396_n6451.n258 0.635332
R6201 a_5396_n6451.n261 a_5396_n6451.n243 0.635332
R6202 a_5396_n6451.n259 a_5396_n6451.n240 0.635332
R6203 a_5396_n6451.n257 a_5396_n6451.n237 0.635332
R6204 a_5396_n6451.n254 a_5396_n6451.n231 0.635332
R6205 a_5396_n6451.n251 a_5396_n6451.n228 0.635332
R6206 a_5396_n6451.n224 a_5396_n6451.n249 0.635332
R6207 a_5396_n6451.n137 a_5396_n6451.n389 0.431935
R6208 a_5396_n6451.n403 a_5396_n6451.n138 0.431935
R6209 a_5396_n6451.n412 a_5396_n6451.n143 0.431935
R6210 a_5396_n6451.n455 a_5396_n6451.n129 0.431935
R6211 a_5396_n6451.n452 a_5396_n6451.n132 0.431935
R6212 a_5396_n6451.n135 a_5396_n6451.n445 0.431935
R6213 a_5396_n6451.n290 a_5396_n6451.n31 0.891677
R6214 a_5396_n6451.n29 a_5396_n6451.n289 0.891677
R6215 a_5396_n6451.n302 a_5396_n6451.n162 0.891728
R6216 a_5396_n6451.n160 a_5396_n6451.n301 0.891728
R6217 a_5396_n6451.n280 a_5396_n6451.n183 0.63266
R6218 a_5396_n6451.n7 a_5396_n6451.n179 0.892822
R6219 a_5396_n6451.n179 a_5396_n6451.n283 0.63266
R6220 a_5396_n6451.n4 a_5396_n6451.n172 1.74336
R6221 a_5396_n6451.n292 a_5396_n6451.n35 0.891677
R6222 a_5396_n6451.n291 a_5396_n6451.n33 0.891677
R6223 a_5396_n6451.n166 a_5396_n6451.n305 0.891728
R6224 a_5396_n6451.n303 a_5396_n6451.n164 0.891728
R6225 a_5396_n6451.n191 a_5396_n6451.n16 0.892462
R6226 a_5396_n6451.n188 a_5396_n6451.n13 0.892822
R6227 a_5396_n6451.n277 a_5396_n6451.n188 0.63266
R6228 a_5396_n6451.n10 a_5396_n6451.n185 1.74336
R6229 a_5396_n6451.n382 a_5396_n6451.n381 0.3605
R6230 a_5396_n6451.n424 a_5396_n6451.n386 0.3605
R6231 a_5396_n6451.n375 a_5396_n6451.n372 0.3605
R6232 a_5396_n6451.n474 a_5396_n6451.n366 0.3605
R6233 a_5396_n6451.n610 a_5396_n6451.n327 0.478684
R6234 a_5396_n6451.n609 a_5396_n6451.n321 0.478684
R6235 a_5396_n6451.n568 a_5396_n6451.n337 0.478684
R6236 a_5396_n6451.n567 a_5396_n6451.n331 0.478684
R6237 a_5396_n6451.n374 a_5396_n6451.n373 0.327481
R6238 a_5396_n6451.n380 a_5396_n6451.n379 0.327481
R6239 a_5396_n6451.n406 a_5396_n6451.n114 0.302474
R6240 a_5396_n6451.n316 a_5396_n6451.n155 0.302474
R6241 a_5396_n6451.n108 a_5396_n6451.n394 0.302474
R6242 a_5396_n6451.n149 a_5396_n6451.n451 0.302474
R6243 a_5396_n6451.n146 a_5396_n6451.n454 0.302474
R6244 a_5396_n6451.n435 a_5396_n6451.n104 0.302474
R6245 a_5396_n6451.n265 a_5396_n6451.n210 0.559597
R6246 a_5396_n6451.n263 a_5396_n6451.n206 0.559597
R6247 a_5396_n6451.n279 a_5396_n6451.n182 0.559597
R6248 a_5396_n6451.n282 a_5396_n6451.n178 0.559597
R6249 a_5396_n6451.n221 a_5396_n6451.n269 0.559597
R6250 a_5396_n6451.n216 a_5396_n6451.n267 0.559597
R6251 a_5396_n6451.n270 a_5396_n6451.n220 0.559597
R6252 a_5396_n6451.n268 a_5396_n6451.n215 0.559597
R6253 a_5396_n6451.n276 a_5396_n6451.n187 0.559597
R6254 a_5396_n6451.n266 a_5396_n6451.n209 0.559597
R6255 a_5396_n6451.n264 a_5396_n6451.n205 0.559597
R6256 a_5396_n6451.n393 a_5396_n6451.n390 0.287375
R6257 a_5396_n6451.n402 a_5396_n6451.n401 0.287375
R6258 a_5396_n6451.n112 a_5396_n6451.n407 0.287375
R6259 a_5396_n6451.n102 a_5396_n6451.n436 0.287375
R6260 a_5396_n6451.n453 a_5396_n6451.n441 0.287375
R6261 a_5396_n6451.n450 a_5396_n6451.n443 0.287375
R6262 a_5396_n6451.n428 a_5396_n6451.n386 0.208099
R6263 a_5396_n6451.n474 a_5396_n6451.n473 0.208099
R6264 a_5396_n6451.n475 a_5396_n6451.n367 0.142605
R6265 a_5396_n6451.n376 a_5396_n6451.n373 0.142605
R6266 a_5396_n6451.n427 a_5396_n6451.n426 0.142605
R6267 a_5396_n6451.n379 a_5396_n6451.n378 0.142605
R6268 a_5396_n6451.n233 a_5396_n6451.n22 0.882326
R6269 a_5396_n6451.n290 a_5396_n6451.n22 1.19478
R6270 a_5396_n6451.n255 a_5396_n6451.n31 1.23157
R6271 a_5396_n6451.n252 a_5396_n6451.n265 3.29744
R6272 a_5396_n6451.n289 a_5396_n6451.n263 0.960161
R6273 a_5396_n6451.n29 a_5396_n6451.n250 1.23157
R6274 a_5396_n6451.n302 a_5396_n6451.n279 0.960134
R6275 a_5396_n6451.n8 a_5396_n6451.n162 1.49213
R6276 a_5396_n6451.n282 a_5396_n6451.n1 3.55769
R6277 a_5396_n6451.n1 a_5396_n6451.n176 0.908313
R6278 a_5396_n6451.n176 a_5396_n6451.n284 0.559957
R6279 a_5396_n6451.n301 a_5396_n6451.n284 0.960134
R6280 a_5396_n6451.n160 a_5396_n6451.n5 1.49213
R6281 a_5396_n6451.n280 a_5396_n6451.n296 0.953788
R6282 a_5396_n6451.n2 a_5396_n6451.n283 3.50093
R6283 a_5396_n6451.n2 a_5396_n6451.n175 0.892822
R6284 a_5396_n6451.n175 a_5396_n6451.n285 0.63302
R6285 a_5396_n6451.n285 a_5396_n6451.n295 0.953788
R6286 a_5396_n6451.n19 a_5396_n6451.n247 0.882326
R6287 a_5396_n6451.n292 a_5396_n6451.n19 1.19478
R6288 a_5396_n6451.n262 a_5396_n6451.n35 1.23157
R6289 a_5396_n6451.n260 a_5396_n6451.n269 3.29744
R6290 a_5396_n6451.n291 a_5396_n6451.n267 0.960161
R6291 a_5396_n6451.n258 a_5396_n6451.n33 1.23157
R6292 a_5396_n6451.n245 a_5396_n6451.n20 0.882326
R6293 a_5396_n6451.n459 a_5396_n6451.n20 1.21084
R6294 a_5396_n6451.n270 a_5396_n6451.n259 3.29744
R6295 a_5396_n6451.n268 a_5396_n6451.n298 0.976221
R6296 a_5396_n6451.n271 a_5396_n6451.n197 0.559957
R6297 a_5396_n6451.n305 a_5396_n6451.n271 0.960134
R6298 a_5396_n6451.n166 a_5396_n6451.n17 1.49213
R6299 a_5396_n6451.n273 a_5396_n6451.n192 0.559957
R6300 a_5396_n6451.n14 a_5396_n6451.n273 3.55805
R6301 a_5396_n6451.n303 a_5396_n6451.n276 0.960134
R6302 a_5396_n6451.n11 a_5396_n6451.n164 1.49213
R6303 a_5396_n6451.n272 a_5396_n6451.n196 0.63302
R6304 a_5396_n6451.n461 a_5396_n6451.n272 0.953788
R6305 a_5396_n6451.n274 a_5396_n6451.n191 0.63302
R6306 a_5396_n6451.n13 a_5396_n6451.n274 3.50129
R6307 a_5396_n6451.n277 a_5396_n6451.n297 0.953788
R6308 a_5396_n6451.n23 a_5396_n6451.n235 0.882326
R6309 a_5396_n6451.n23 a_5396_n6451.n299 1.21084
R6310 a_5396_n6451.n266 a_5396_n6451.n251 3.29744
R6311 a_5396_n6451.n264 a_5396_n6451.n464 0.976221
R6312 a_5396_n6451.n307 a_5396_n6451.n391 1.12843
R6313 a_5396_n6451.n393 a_5396_n6451.n153 0.209185
R6314 a_5396_n6451.n110 a_5396_n6451.n390 0.209185
R6315 a_5396_n6451.n377 a_5396_n6451.n110 2.25894
R6316 a_5396_n6451.n123 a_5396_n6451.n389 0.209185
R6317 a_5396_n6451.n399 a_5396_n6451.n137 0.209185
R6318 a_5396_n6451.n401 a_5396_n6451.n154 0.209185
R6319 a_5396_n6451.n402 a_5396_n6451.n318 0.208307
R6320 a_5396_n6451.n312 a_5396_n6451.n318 3.16466
R6321 a_5396_n6451.n403 a_5396_n6451.n312 0.208324
R6322 a_5396_n6451.n405 a_5396_n6451.n138 0.209185
R6323 a_5396_n6451.n407 a_5396_n6451.n158 0.209185
R6324 a_5396_n6451.n113 a_5396_n6451.n112 0.209185
R6325 a_5396_n6451.n113 a_5396_n6451.n111 2.25894
R6326 a_5396_n6451.n412 a_5396_n6451.n126 0.209185
R6327 a_5396_n6451.n143 a_5396_n6451.n411 0.209185
R6328 a_5396_n6451.n382 a_5396_n6451.n51 0.209185
R6329 a_5396_n6451.n45 a_5396_n6451.n51 0.429685
R6330 a_5396_n6451.n46 a_5396_n6451.n45 0.209185
R6331 a_5396_n6451.n46 a_5396_n6451.n44 2.23644
R6332 a_5396_n6451.n432 a_5396_n6451.n59 0.209185
R6333 a_5396_n6451.n430 a_5396_n6451.n59 0.429685
R6334 a_5396_n6451.n430 a_5396_n6451.n55 0.209185
R6335 a_5396_n6451.n55 a_5396_n6451.n54 0.429685
R6336 a_5396_n6451.n54 a_5396_n6451.n53 0.209185
R6337 a_5396_n6451.n53 a_5396_n6451.n37 0.564455
R6338 a_5396_n6451.n37 a_5396_n6451.n428 3.17649
R6339 a_5396_n6451.n424 a_5396_n6451.n65 0.209185
R6340 a_5396_n6451.n65 a_5396_n6451.n387 0.429685
R6341 a_5396_n6451.n63 a_5396_n6451.n387 0.209185
R6342 a_5396_n6451.n63 a_5396_n6451.n388 0.429685
R6343 a_5396_n6451.n61 a_5396_n6451.n388 0.209185
R6344 a_5396_n6451.n61 a_5396_n6451.n414 2.23644
R6345 a_5396_n6451.n417 a_5396_n6451.n69 0.209185
R6346 a_5396_n6451.n69 a_5396_n6451.n415 0.429685
R6347 a_5396_n6451.n67 a_5396_n6451.n415 0.209185
R6348 a_5396_n6451.n67 a_5396_n6451.n38 1.26163
R6349 a_5396_n6451.n434 a_5396_n6451.n308 1.12843
R6350 a_5396_n6451.n436 a_5396_n6451.n145 0.209185
R6351 a_5396_n6451.n103 a_5396_n6451.n102 0.209185
R6352 a_5396_n6451.n103 a_5396_n6451.n101 2.25894
R6353 a_5396_n6451.n455 a_5396_n6451.n118 0.209185
R6354 a_5396_n6451.n129 a_5396_n6451.n440 0.209185
R6355 a_5396_n6451.n148 a_5396_n6451.n441 0.209185
R6356 a_5396_n6451.n453 a_5396_n6451.n320 0.208307
R6357 a_5396_n6451.n320 a_5396_n6451.n315 3.16466
R6358 a_5396_n6451.n452 a_5396_n6451.n315 0.208324
R6359 a_5396_n6451.n132 a_5396_n6451.n442 0.209185
R6360 a_5396_n6451.n151 a_5396_n6451.n443 0.209185
R6361 a_5396_n6451.n450 a_5396_n6451.n107 0.209185
R6362 a_5396_n6451.n107 a_5396_n6451.n444 2.25894
R6363 a_5396_n6451.n121 a_5396_n6451.n445 0.209185
R6364 a_5396_n6451.n135 a_5396_n6451.n446 0.209185
R6365 a_5396_n6451.n75 a_5396_n6451.n372 0.209185
R6366 a_5396_n6451.n371 a_5396_n6451.n75 0.429685
R6367 a_5396_n6451.n72 a_5396_n6451.n371 0.209185
R6368 a_5396_n6451.n469 a_5396_n6451.n72 2.23644
R6369 a_5396_n6451.n84 a_5396_n6451.n370 0.209185
R6370 a_5396_n6451.n369 a_5396_n6451.n84 0.429685
R6371 a_5396_n6451.n81 a_5396_n6451.n369 0.209185
R6372 a_5396_n6451.n368 a_5396_n6451.n81 0.429685
R6373 a_5396_n6451.n78 a_5396_n6451.n368 0.209185
R6374 a_5396_n6451.n41 a_5396_n6451.n78 0.564455
R6375 a_5396_n6451.n473 a_5396_n6451.n41 3.17649
R6376 a_5396_n6451.n95 a_5396_n6451.n366 0.209185
R6377 a_5396_n6451.n476 a_5396_n6451.n95 0.429685
R6378 a_5396_n6451.n476 a_5396_n6451.n92 0.209185
R6379 a_5396_n6451.n86 a_5396_n6451.n92 0.429685
R6380 a_5396_n6451.n87 a_5396_n6451.n86 0.209185
R6381 a_5396_n6451.n87 a_5396_n6451.n85 2.23644
R6382 a_5396_n6451.n482 a_5396_n6451.n100 0.209185
R6383 a_5396_n6451.n480 a_5396_n6451.n100 0.429685
R6384 a_5396_n6451.n480 a_5396_n6451.n96 0.209185
R6385 a_5396_n6451.n96 a_5396_n6451.n43 1.26163
R6386 a_5396_n6451.n329 a_5396_n6451.n330 1.27228
R6387 a_5396_n6451.n328 a_5396_n6451.n329 2.51878
R6388 a_5396_n6451.n610 a_5396_n6451.n328 0.794091
R6389 a_5396_n6451.n326 a_5396_n6451.n327 1.27228
R6390 a_5396_n6451.n325 a_5396_n6451.n326 2.60203
R6391 a_5396_n6451.n324 a_5396_n6451.n325 1.27228
R6392 a_5396_n6451.n323 a_5396_n6451.n324 1.27228
R6393 a_5396_n6451.n322 a_5396_n6451.n323 2.51878
R6394 a_5396_n6451.n609 a_5396_n6451.n322 0.794091
R6395 a_5396_n6451.t39 a_5396_n6451.n321 6.77266
R6396 a_5396_n6451.n339 a_5396_n6451.n340 1.27228
R6397 a_5396_n6451.n338 a_5396_n6451.n339 2.51878
R6398 a_5396_n6451.n568 a_5396_n6451.n338 0.794091
R6399 a_5396_n6451.n336 a_5396_n6451.n337 1.27228
R6400 a_5396_n6451.n335 a_5396_n6451.n336 2.60203
R6401 a_5396_n6451.n334 a_5396_n6451.n335 1.27228
R6402 a_5396_n6451.n333 a_5396_n6451.n334 1.27228
R6403 a_5396_n6451.n332 a_5396_n6451.n333 2.51878
R6404 a_5396_n6451.n567 a_5396_n6451.n332 0.794091
R6405 a_5396_n6451.t20 a_5396_n6451.n331 6.77266
R6406 a_5396_n6451.n531 a_5396_n6451.n341 3.17898
R6407 a_5396_n6451.n40 a_5396_n6451.n77 0.531026
R6408 a_5396_n6451.n52 a_5396_n6451.n36 0.531026
R6409 a_5396_n6451.n34 a_5396_n6451.n202 0.386311
R6410 a_5396_n6451.n32 a_5396_n6451.n201 0.386311
R6411 a_5396_n6451.n30 a_5396_n6451.n200 0.386311
R6412 a_5396_n6451.n288 a_5396_n6451.n28 0.386311
R6413 a_5396_n6451.n304 a_5396_n6451.n165 0.364343
R6414 a_5396_n6451.n163 a_5396_n6451.n287 0.364343
R6415 a_5396_n6451.n161 a_5396_n6451.n286 0.364343
R6416 a_5396_n6451.n300 a_5396_n6451.n159 0.364343
R6417 a_5396_n6451.n190 a_5396_n6451.n15 0.354735
R6418 a_5396_n6451.n186 a_5396_n6451.n12 0.354735
R6419 a_5396_n6451.n184 a_5396_n6451.n9 0.354735
R6420 a_5396_n6451.n177 a_5396_n6451.n6 0.354735
R6421 a_5396_n6451.n3 a_5396_n6451.n171 0.354735
R6422 a_5396_n6451.n0 a_5396_n6451.n174 0.354735
R6423 a_5396_n6451.n21 a_5396_n6451.n211 0.347689
R6424 a_5396_n6451.n18 a_5396_n6451.n222 0.347689
R6425 a_5396_n6451.n406 a_5396_n6451.n157 0.294184
R6426 a_5396_n6451.n156 a_5396_n6451.n155 0.294184
R6427 a_5396_n6451.n394 a_5396_n6451.n152 0.294184
R6428 a_5396_n6451.n150 a_5396_n6451.n149 0.294184
R6429 a_5396_n6451.n147 a_5396_n6451.n146 0.294184
R6430 a_5396_n6451.n435 a_5396_n6451.n144 0.294184
R6431 a_5396_n6451.n142 a_5396_n6451.n141 0.294184
R6432 a_5396_n6451.n140 a_5396_n6451.n139 0.294184
R6433 a_5396_n6451.n400 a_5396_n6451.n136 0.294184
R6434 a_5396_n6451.n134 a_5396_n6451.n133 0.294184
R6435 a_5396_n6451.n131 a_5396_n6451.n130 0.294184
R6436 a_5396_n6451.n128 a_5396_n6451.n127 0.294184
R6437 a_5396_n6451.n125 a_5396_n6451.n124 0.294184
R6438 a_5396_n6451.n398 a_5396_n6451.n122 0.294184
R6439 a_5396_n6451.n120 a_5396_n6451.n119 0.294184
R6440 a_5396_n6451.n117 a_5396_n6451.n116 0.294184
R6441 a_5396_n6451.n115 a_5396_n6451.n114 0.294184
R6442 a_5396_n6451.n109 a_5396_n6451.n108 0.294184
R6443 a_5396_n6451.n451 a_5396_n6451.n106 0.294184
R6444 a_5396_n6451.n105 a_5396_n6451.n104 0.294184
R6445 a_5396_n6451.n481 a_5396_n6451.n99 0.294184
R6446 a_5396_n6451.n98 a_5396_n6451.n97 0.294184
R6447 a_5396_n6451.n94 a_5396_n6451.n93 0.294184
R6448 a_5396_n6451.n91 a_5396_n6451.n90 0.294184
R6449 a_5396_n6451.n89 a_5396_n6451.n88 0.294184
R6450 a_5396_n6451.n83 a_5396_n6451.n82 0.294184
R6451 a_5396_n6451.n80 a_5396_n6451.n79 0.294184
R6452 a_5396_n6451.n77 a_5396_n6451.n76 0.294184
R6453 a_5396_n6451.n74 a_5396_n6451.n73 0.294184
R6454 a_5396_n6451.n71 a_5396_n6451.n70 0.294184
R6455 a_5396_n6451.n418 a_5396_n6451.n68 0.294184
R6456 a_5396_n6451.n416 a_5396_n6451.n66 0.294184
R6457 a_5396_n6451.n425 a_5396_n6451.n64 0.294184
R6458 a_5396_n6451.n423 a_5396_n6451.n62 0.294184
R6459 a_5396_n6451.n422 a_5396_n6451.n60 0.294184
R6460 a_5396_n6451.n431 a_5396_n6451.n58 0.294184
R6461 a_5396_n6451.n57 a_5396_n6451.n56 0.294184
R6462 a_5396_n6451.n429 a_5396_n6451.n52 0.294184
R6463 a_5396_n6451.n50 a_5396_n6451.n49 0.294184
R6464 a_5396_n6451.n48 a_5396_n6451.n47 0.294184
R6465 a_5396_n6451.n195 a_5396_n6451.n194 0.255447
R6466 a_5396_n6451.n190 a_5396_n6451.n189 0.255447
R6467 a_5396_n6451.n275 a_5396_n6451.n186 0.255447
R6468 a_5396_n6451.n278 a_5396_n6451.n181 0.255447
R6469 a_5396_n6451.n281 a_5396_n6451.n177 0.255447
R6470 a_5396_n6451.n174 a_5396_n6451.n173 0.255447
R6471 a_5396_n6451.n219 a_5396_n6451.n218 0.241034
R6472 a_5396_n6451.n214 a_5396_n6451.n213 0.241034
R6473 a_5396_n6451.n208 a_5396_n6451.n207 0.241034
R6474 a_5396_n6451.n204 a_5396_n6451.n203 0.241034
R6475 a_5396_n6451.n219 a_5396_n6451.n217 0.186585
R6476 a_5396_n6451.n214 a_5396_n6451.n212 0.186585
R6477 a_5396_n6451.n236 a_5396_n6451.n24 0.186585
R6478 a_5396_n6451.n230 a_5396_n6451.n208 0.186585
R6479 a_5396_n6451.n227 a_5396_n6451.n204 0.186585
R6480 a_5396_n6451.n223 a_5396_n6451.n26 0.186585
R6481 a_5396_n6451.n217 a_5396_n6451.n242 0.183062
R6482 a_5396_n6451.n212 a_5396_n6451.n239 0.183062
R6483 a_5396_n6451.n256 a_5396_n6451.n236 0.183062
R6484 a_5396_n6451.n253 a_5396_n6451.n230 0.183062
R6485 a_5396_n6451.n227 a_5396_n6451.n226 0.183062
R6486 a_5396_n6451.n248 a_5396_n6451.n223 0.183062
R6487 a_5396_n6451.n222 a_5396_n6451.n246 0.183062
R6488 a_5396_n6451.n211 a_5396_n6451.n234 0.183062
R6489 a_5396_n6451.n195 a_5396_n6451.n193 0.182422
R6490 a_5396_n6451.n181 a_5396_n6451.n180 0.182422
R6491 a_5396_n6451.n310 a_5396_n6451.n309 0.1805
R6492 a_5396_n6451.n392 a_5396_n6451.n306 0.1805
R6493 a_5396_n6451.n314 a_5396_n6451.n313 0.178132
R6494 a_5396_n6451.n404 a_5396_n6451.n311 0.178132
R6495 a_5396_n6451.n454 a_5396_n6451.n319 0.175763
R6496 a_5396_n6451.n317 a_5396_n6451.n316 0.175763
R6497 a_5396_8177.n90 a_5396_8177.n89 7.22198
R6498 a_5396_8177.n262 a_5396_8177.n261 7.22198
R6499 a_5396_8177.n50 a_5396_8177.n47 6.77653
R6500 a_5396_8177.n43 a_5396_8177.n40 6.77653
R6501 a_5396_8177.n56 a_5396_8177.t41 6.7761
R6502 a_5396_8177.n280 a_5396_8177.t80 6.7761
R6503 a_5396_8177.n8 a_5396_8177.n92 6.77231
R6504 a_5396_8177.n18 a_5396_8177.n102 6.77231
R6505 a_5396_8177.n221 a_5396_8177.n220 6.50088
R6506 a_5396_8177.n174 a_5396_8177.n168 6.50088
R6507 a_5396_8177.n60 a_5396_8177.t21 5.50607
R6508 a_5396_8177.n51 a_5396_8177.t28 5.50607
R6509 a_5396_8177.n275 a_5396_8177.t56 5.50607
R6510 a_5396_8177.n44 a_5396_8177.t66 5.50607
R6511 a_5396_8177.n59 a_5396_8177.n58 5.50475
R6512 a_5396_8177.n65 a_5396_8177.n64 5.50475
R6513 a_5396_8177.n66 a_5396_8177.t54 5.50475
R6514 a_5396_8177.n53 a_5396_8177.n52 5.50475
R6515 a_5396_8177.n277 a_5396_8177.n276 5.50475
R6516 a_5396_8177.n271 a_5396_8177.n270 5.50475
R6517 a_5396_8177.n269 a_5396_8177.t4 5.50475
R6518 a_5396_8177.n46 a_5396_8177.n45 5.50475
R6519 a_5396_8177.n119 a_5396_8177.n116 4.92758
R6520 a_5396_8177.n182 a_5396_8177.n179 4.92758
R6521 a_5396_8177.n25 a_5396_8177.n128 4.92217
R6522 a_5396_8177.n32 a_5396_8177.n151 4.92217
R6523 a_5396_8177.n19 a_5396_8177.n142 3.65107
R6524 a_5396_8177.n20 a_5396_8177.n140 3.65107
R6525 a_5396_8177.n21 a_5396_8177.n138 3.65107
R6526 a_5396_8177.n22 a_5396_8177.n136 3.65107
R6527 a_5396_8177.n134 a_5396_8177.n23 3.65107
R6528 a_5396_8177.n132 a_5396_8177.n24 3.65107
R6529 a_5396_8177.n130 a_5396_8177.n25 3.65107
R6530 a_5396_8177.n26 a_5396_8177.n165 3.65107
R6531 a_5396_8177.n27 a_5396_8177.n163 3.65107
R6532 a_5396_8177.n28 a_5396_8177.n161 3.65107
R6533 a_5396_8177.n29 a_5396_8177.n159 3.65107
R6534 a_5396_8177.n157 a_5396_8177.n30 3.65107
R6535 a_5396_8177.n155 a_5396_8177.n31 3.65107
R6536 a_5396_8177.n153 a_5396_8177.n32 3.65107
R6537 a_5396_8177.n33 a_5396_8177.n285 4.0312
R6538 a_5396_8177.n0 a_5396_8177.n37 4.0312
R6539 a_5396_8177.n1 a_5396_8177.n35 5.5012
R6540 a_5396_8177.n2 a_5396_8177.t32 5.5012
R6541 a_5396_8177.n3 a_5396_8177.n98 5.5012
R6542 a_5396_8177.n4 a_5396_8177.t67 5.5012
R6543 a_5396_8177.n5 a_5396_8177.n97 4.0312
R6544 a_5396_8177.n95 a_5396_8177.n6 5.5012
R6545 a_5396_8177.t39 a_5396_8177.n7 5.5012
R6546 a_5396_8177.n94 a_5396_8177.n8 4.0312
R6547 a_5396_8177.n9 a_5396_8177.n113 4.0312
R6548 a_5396_8177.n10 a_5396_8177.n111 5.5012
R6549 a_5396_8177.n11 a_5396_8177.t79 5.5012
R6550 a_5396_8177.n12 a_5396_8177.n110 4.0312
R6551 a_5396_8177.n13 a_5396_8177.n108 5.5012
R6552 a_5396_8177.n14 a_5396_8177.t37 5.5012
R6553 a_5396_8177.n15 a_5396_8177.n107 4.0312
R6554 a_5396_8177.n105 a_5396_8177.n16 5.5012
R6555 a_5396_8177.t42 a_5396_8177.n17 5.5012
R6556 a_5396_8177.n104 a_5396_8177.n18 4.0312
R6557 a_5396_8177.n88 a_5396_8177.n87 4.24002
R6558 a_5396_8177.n73 a_5396_8177.n72 4.24002
R6559 a_5396_8177.n260 a_5396_8177.n259 4.24002
R6560 a_5396_8177.n245 a_5396_8177.n244 4.24002
R6561 a_5396_8177.n175 a_5396_8177.t134 4.06712
R6562 a_5396_8177.n148 a_5396_8177.t143 4.06712
R6563 a_5396_8177.n213 a_5396_8177.t124 4.06712
R6564 a_5396_8177.n211 a_5396_8177.t166 4.06712
R6565 a_5396_8177.n56 a_5396_8177.n55 4.03475
R6566 a_5396_8177.n63 a_5396_8177.n62 4.03475
R6567 a_5396_8177.n69 a_5396_8177.n68 4.03475
R6568 a_5396_8177.n50 a_5396_8177.n49 4.03475
R6569 a_5396_8177.n280 a_5396_8177.n279 4.03475
R6570 a_5396_8177.n274 a_5396_8177.n273 4.03475
R6571 a_5396_8177.n268 a_5396_8177.n267 4.03475
R6572 a_5396_8177.n43 a_5396_8177.n42 4.03475
R6573 a_5396_8177.n238 a_5396_8177.n101 3.97307
R6574 a_5396_8177.n214 a_5396_8177.n114 3.96014
R6575 a_5396_8177.n177 a_5396_8177.n176 3.96014
R6576 a_5396_8177.n175 a_5396_8177.t133 3.86107
R6577 a_5396_8177.n148 a_5396_8177.t142 3.86107
R6578 a_5396_8177.n213 a_5396_8177.t125 3.86107
R6579 a_5396_8177.n211 a_5396_8177.t168 3.86107
R6580 a_5396_8177.n122 a_5396_8177.n119 3.79678
R6581 a_5396_8177.n233 a_5396_8177.n230 3.79678
R6582 a_5396_8177.n185 a_5396_8177.n182 3.79678
R6583 a_5396_8177.n198 a_5396_8177.n195 3.79678
R6584 a_5396_8177.n88 a_5396_8177.n86 3.68818
R6585 a_5396_8177.n73 a_5396_8177.n71 3.68818
R6586 a_5396_8177.n260 a_5396_8177.n258 3.68818
R6587 a_5396_8177.n245 a_5396_8177.n243 3.68818
R6588 a_5396_8177.n236 a_5396_8177.n235 3.65581
R6589 a_5396_8177.n233 a_5396_8177.n232 3.65581
R6590 a_5396_8177.n230 a_5396_8177.n229 3.65581
R6591 a_5396_8177.n227 a_5396_8177.n226 3.65581
R6592 a_5396_8177.n125 a_5396_8177.n124 3.65581
R6593 a_5396_8177.n122 a_5396_8177.n121 3.65581
R6594 a_5396_8177.n119 a_5396_8177.n118 3.65581
R6595 a_5396_8177.n201 a_5396_8177.n200 3.65581
R6596 a_5396_8177.n198 a_5396_8177.n197 3.65581
R6597 a_5396_8177.n195 a_5396_8177.n194 3.65581
R6598 a_5396_8177.n192 a_5396_8177.n191 3.65581
R6599 a_5396_8177.n188 a_5396_8177.n187 3.65581
R6600 a_5396_8177.n185 a_5396_8177.n184 3.65581
R6601 a_5396_8177.n182 a_5396_8177.n181 3.65581
R6602 a_5396_8177.n227 a_5396_8177.n224 3.64443
R6603 a_5396_8177.n192 a_5396_8177.n189 3.64443
R6604 a_5396_8177.n204 a_5396_8177.n22 3.64223
R6605 a_5396_8177.n166 a_5396_8177.n29 3.64223
R6606 a_5396_8177.n85 a_5396_8177.n38 3.23904
R6607 a_5396_8177.n257 a_5396_8177.n39 3.23904
R6608 a_5396_8177.n84 a_5396_8177.n83 2.77002
R6609 a_5396_8177.n78 a_5396_8177.n77 2.77002
R6610 a_5396_8177.n256 a_5396_8177.n255 2.77002
R6611 a_5396_8177.n250 a_5396_8177.n249 2.77002
R6612 a_5396_8177.n79 a_5396_8177.n73 2.73714
R6613 a_5396_8177.n251 a_5396_8177.n245 2.73714
R6614 a_5396_8177.n212 a_5396_8177.n210 2.73714
R6615 a_5396_8177.n149 a_5396_8177.n147 2.73714
R6616 a_5396_8177.n66 a_5396_8177.n65 2.60203
R6617 a_5396_8177.n271 a_5396_8177.n269 2.60203
R6618 a_5396_8177.n173 a_5396_8177.n170 2.59712
R6619 a_5396_8177.n147 a_5396_8177.n144 2.59712
R6620 a_5396_8177.n219 a_5396_8177.n216 2.59712
R6621 a_5396_8177.n210 a_5396_8177.n207 2.59712
R6622 a_5396_8177.n53 a_5396_8177.n51 2.52436
R6623 a_5396_8177.n60 a_5396_8177.n59 2.52436
R6624 a_5396_8177.n46 a_5396_8177.n44 2.52436
R6625 a_5396_8177.n277 a_5396_8177.n275 2.52436
R6626 a_5396_8177.n221 a_5396_8177.n212 2.46014
R6627 a_5396_8177.n168 a_5396_8177.n149 2.46014
R6628 a_5396_8177.n173 a_5396_8177.n172 2.39107
R6629 a_5396_8177.n147 a_5396_8177.n146 2.39107
R6630 a_5396_8177.n219 a_5396_8177.n218 2.39107
R6631 a_5396_8177.n210 a_5396_8177.n209 2.39107
R6632 a_5396_8177.n84 a_5396_8177.n81 2.21818
R6633 a_5396_8177.n78 a_5396_8177.n75 2.21818
R6634 a_5396_8177.n256 a_5396_8177.n253 2.21818
R6635 a_5396_8177.n250 a_5396_8177.n247 2.21818
R6636 a_5396_8177.n91 a_5396_8177.n70 2.13841
R6637 a_5396_8177.n57 a_5396_8177.n38 2.13841
R6638 a_5396_8177.n167 a_5396_8177.n166 2.0852
R6639 a_5396_8177.n238 a_5396_8177.n237 2.02864
R6640 a_5396_8177.n242 a_5396_8177.n101 1.76168
R6641 a_5396_8177.n90 a_5396_8177.n79 1.73904
R6642 a_5396_8177.n262 a_5396_8177.n251 1.73904
R6643 a_5396_8177.n237 a_5396_8177.n236 1.73609
R6644 a_5396_8177.n202 a_5396_8177.n201 1.73609
R6645 a_5396_8177.n242 a_5396_8177.n241 1.5005
R6646 a_5396_8177.n263 a_5396_8177.n262 1.5005
R6647 a_5396_8177.n265 a_5396_8177.n264 1.5005
R6648 a_5396_8177.n91 a_5396_8177.n90 1.5005
R6649 a_5396_8177.n222 a_5396_8177.n221 1.5005
R6650 a_5396_8177.n189 a_5396_8177.n126 1.5005
R6651 a_5396_8177.n205 a_5396_8177.n204 1.5005
R6652 a_5396_8177.n224 a_5396_8177.n223 1.5005
R6653 a_5396_8177.n168 a_5396_8177.n167 1.5005
R6654 a_5396_8177.n240 a_5396_8177.n239 1.5005
R6655 a_5396_8177.n282 a_5396_8177.n281 1.5005
R6656 a_5396_8177.n284 a_5396_8177.n283 1.5005
R6657 a_5396_8177.n100 a_5396_8177.n99 1.5005
R6658 a_5396_8177.n37 a_5396_8177.t44 1.4705
R6659 a_5396_8177.n37 a_5396_8177.n36 1.4705
R6660 a_5396_8177.n97 a_5396_8177.t35 1.4705
R6661 a_5396_8177.n97 a_5396_8177.n96 1.4705
R6662 a_5396_8177.n94 a_5396_8177.t81 1.4705
R6663 a_5396_8177.n94 a_5396_8177.n93 1.4705
R6664 a_5396_8177.n55 a_5396_8177.t33 1.4705
R6665 a_5396_8177.n55 a_5396_8177.n54 1.4705
R6666 a_5396_8177.n62 a_5396_8177.t76 1.4705
R6667 a_5396_8177.n62 a_5396_8177.n61 1.4705
R6668 a_5396_8177.n68 a_5396_8177.t22 1.4705
R6669 a_5396_8177.n68 a_5396_8177.n67 1.4705
R6670 a_5396_8177.n49 a_5396_8177.t68 1.4705
R6671 a_5396_8177.n49 a_5396_8177.n48 1.4705
R6672 a_5396_8177.n81 a_5396_8177.t72 1.4705
R6673 a_5396_8177.n81 a_5396_8177.n80 1.4705
R6674 a_5396_8177.n83 a_5396_8177.t74 1.4705
R6675 a_5396_8177.n83 a_5396_8177.n82 1.4705
R6676 a_5396_8177.n75 a_5396_8177.t83 1.4705
R6677 a_5396_8177.n75 a_5396_8177.n74 1.4705
R6678 a_5396_8177.n77 a_5396_8177.t1 1.4705
R6679 a_5396_8177.n77 a_5396_8177.n76 1.4705
R6680 a_5396_8177.n279 a_5396_8177.t71 1.4705
R6681 a_5396_8177.n279 a_5396_8177.n278 1.4705
R6682 a_5396_8177.n273 a_5396_8177.t26 1.4705
R6683 a_5396_8177.n273 a_5396_8177.n272 1.4705
R6684 a_5396_8177.n267 a_5396_8177.t59 1.4705
R6685 a_5396_8177.n267 a_5396_8177.n266 1.4705
R6686 a_5396_8177.n42 a_5396_8177.t18 1.4705
R6687 a_5396_8177.n42 a_5396_8177.n41 1.4705
R6688 a_5396_8177.n253 a_5396_8177.t19 1.4705
R6689 a_5396_8177.n253 a_5396_8177.n252 1.4705
R6690 a_5396_8177.n255 a_5396_8177.t70 1.4705
R6691 a_5396_8177.n255 a_5396_8177.n254 1.4705
R6692 a_5396_8177.n247 a_5396_8177.t31 1.4705
R6693 a_5396_8177.n247 a_5396_8177.n246 1.4705
R6694 a_5396_8177.n249 a_5396_8177.t27 1.4705
R6695 a_5396_8177.n249 a_5396_8177.n248 1.4705
R6696 a_5396_8177.n113 a_5396_8177.t36 1.4705
R6697 a_5396_8177.n113 a_5396_8177.n112 1.4705
R6698 a_5396_8177.n110 a_5396_8177.t57 1.4705
R6699 a_5396_8177.n110 a_5396_8177.n109 1.4705
R6700 a_5396_8177.n107 a_5396_8177.t16 1.4705
R6701 a_5396_8177.n107 a_5396_8177.n106 1.4705
R6702 a_5396_8177.n104 a_5396_8177.t8 1.4705
R6703 a_5396_8177.n104 a_5396_8177.n103 1.4705
R6704 a_5396_8177.n170 a_5396_8177.t95 1.4705
R6705 a_5396_8177.n170 a_5396_8177.n169 1.4705
R6706 a_5396_8177.n172 a_5396_8177.t93 1.4705
R6707 a_5396_8177.n172 a_5396_8177.n171 1.4705
R6708 a_5396_8177.n144 a_5396_8177.t106 1.4705
R6709 a_5396_8177.n144 a_5396_8177.n143 1.4705
R6710 a_5396_8177.n146 a_5396_8177.t105 1.4705
R6711 a_5396_8177.n146 a_5396_8177.n145 1.4705
R6712 a_5396_8177.n235 a_5396_8177.t103 1.4705
R6713 a_5396_8177.n235 a_5396_8177.n234 1.4705
R6714 a_5396_8177.n232 a_5396_8177.t169 1.4705
R6715 a_5396_8177.n232 a_5396_8177.n231 1.4705
R6716 a_5396_8177.n229 a_5396_8177.t156 1.4705
R6717 a_5396_8177.n229 a_5396_8177.n228 1.4705
R6718 a_5396_8177.n226 a_5396_8177.t136 1.4705
R6719 a_5396_8177.n226 a_5396_8177.n225 1.4705
R6720 a_5396_8177.n124 a_5396_8177.t172 1.4705
R6721 a_5396_8177.n124 a_5396_8177.n123 1.4705
R6722 a_5396_8177.n121 a_5396_8177.t150 1.4705
R6723 a_5396_8177.n121 a_5396_8177.n120 1.4705
R6724 a_5396_8177.n118 a_5396_8177.t121 1.4705
R6725 a_5396_8177.n118 a_5396_8177.n117 1.4705
R6726 a_5396_8177.n116 a_5396_8177.t88 1.4705
R6727 a_5396_8177.n116 a_5396_8177.n115 1.4705
R6728 a_5396_8177.n142 a_5396_8177.t158 1.4705
R6729 a_5396_8177.n142 a_5396_8177.n141 1.4705
R6730 a_5396_8177.n140 a_5396_8177.t160 1.4705
R6731 a_5396_8177.n140 a_5396_8177.n139 1.4705
R6732 a_5396_8177.n138 a_5396_8177.t115 1.4705
R6733 a_5396_8177.n138 a_5396_8177.n137 1.4705
R6734 a_5396_8177.n136 a_5396_8177.t137 1.4705
R6735 a_5396_8177.n136 a_5396_8177.n135 1.4705
R6736 a_5396_8177.n134 a_5396_8177.t94 1.4705
R6737 a_5396_8177.n134 a_5396_8177.n133 1.4705
R6738 a_5396_8177.n132 a_5396_8177.t116 1.4705
R6739 a_5396_8177.n132 a_5396_8177.n131 1.4705
R6740 a_5396_8177.n130 a_5396_8177.t148 1.4705
R6741 a_5396_8177.n130 a_5396_8177.n129 1.4705
R6742 a_5396_8177.n128 a_5396_8177.t175 1.4705
R6743 a_5396_8177.n128 a_5396_8177.n127 1.4705
R6744 a_5396_8177.n200 a_5396_8177.t165 1.4705
R6745 a_5396_8177.n200 a_5396_8177.n199 1.4705
R6746 a_5396_8177.n197 a_5396_8177.t130 1.4705
R6747 a_5396_8177.n197 a_5396_8177.n196 1.4705
R6748 a_5396_8177.n194 a_5396_8177.t107 1.4705
R6749 a_5396_8177.n194 a_5396_8177.n193 1.4705
R6750 a_5396_8177.n191 a_5396_8177.t159 1.4705
R6751 a_5396_8177.n191 a_5396_8177.n190 1.4705
R6752 a_5396_8177.n187 a_5396_8177.t151 1.4705
R6753 a_5396_8177.n187 a_5396_8177.n186 1.4705
R6754 a_5396_8177.n184 a_5396_8177.t120 1.4705
R6755 a_5396_8177.n184 a_5396_8177.n183 1.4705
R6756 a_5396_8177.n181 a_5396_8177.t117 1.4705
R6757 a_5396_8177.n181 a_5396_8177.n180 1.4705
R6758 a_5396_8177.n179 a_5396_8177.t155 1.4705
R6759 a_5396_8177.n179 a_5396_8177.n178 1.4705
R6760 a_5396_8177.n165 a_5396_8177.t96 1.4705
R6761 a_5396_8177.n165 a_5396_8177.n164 1.4705
R6762 a_5396_8177.n163 a_5396_8177.t140 1.4705
R6763 a_5396_8177.n163 a_5396_8177.n162 1.4705
R6764 a_5396_8177.n161 a_5396_8177.t122 1.4705
R6765 a_5396_8177.n161 a_5396_8177.n160 1.4705
R6766 a_5396_8177.n159 a_5396_8177.t91 1.4705
R6767 a_5396_8177.n159 a_5396_8177.n158 1.4705
R6768 a_5396_8177.n157 a_5396_8177.t163 1.4705
R6769 a_5396_8177.n157 a_5396_8177.n156 1.4705
R6770 a_5396_8177.n155 a_5396_8177.t135 1.4705
R6771 a_5396_8177.n155 a_5396_8177.n154 1.4705
R6772 a_5396_8177.n153 a_5396_8177.t131 1.4705
R6773 a_5396_8177.n153 a_5396_8177.n152 1.4705
R6774 a_5396_8177.n151 a_5396_8177.t167 1.4705
R6775 a_5396_8177.n151 a_5396_8177.n150 1.4705
R6776 a_5396_8177.n216 a_5396_8177.t99 1.4705
R6777 a_5396_8177.n216 a_5396_8177.n215 1.4705
R6778 a_5396_8177.n218 a_5396_8177.t102 1.4705
R6779 a_5396_8177.n218 a_5396_8177.n217 1.4705
R6780 a_5396_8177.n207 a_5396_8177.t145 1.4705
R6781 a_5396_8177.n207 a_5396_8177.n206 1.4705
R6782 a_5396_8177.n209 a_5396_8177.t146 1.4705
R6783 a_5396_8177.n209 a_5396_8177.n208 1.4705
R6784 a_5396_8177.t87 a_5396_8177.n285 1.4705
R6785 a_5396_8177.n285 a_5396_8177.n34 1.4705
R6786 a_5396_8177.n85 a_5396_8177.n84 1.46537
R6787 a_5396_8177.n89 a_5396_8177.n88 1.46537
R6788 a_5396_8177.n79 a_5396_8177.n78 1.46537
R6789 a_5396_8177.n257 a_5396_8177.n256 1.46537
R6790 a_5396_8177.n261 a_5396_8177.n260 1.46537
R6791 a_5396_8177.n251 a_5396_8177.n250 1.46537
R6792 a_5396_8177.n176 a_5396_8177.n175 1.46537
R6793 a_5396_8177.n174 a_5396_8177.n173 1.46537
R6794 a_5396_8177.n149 a_5396_8177.n148 1.46537
R6795 a_5396_8177.n214 a_5396_8177.n213 1.46537
R6796 a_5396_8177.n220 a_5396_8177.n219 1.46537
R6797 a_5396_8177.n212 a_5396_8177.n211 1.46537
R6798 a_5396_8177.n223 a_5396_8177.n101 1.42428
R6799 a_5396_8177.n69 a_5396_8177.n66 1.27228
R6800 a_5396_8177.n65 a_5396_8177.n63 1.27228
R6801 a_5396_8177.n89 a_5396_8177.n85 1.27228
R6802 a_5396_8177.n269 a_5396_8177.n268 1.27228
R6803 a_5396_8177.n274 a_5396_8177.n271 1.27228
R6804 a_5396_8177.n261 a_5396_8177.n257 1.27228
R6805 a_5396_8177.n125 a_5396_8177.n122 1.27228
R6806 a_5396_8177.n230 a_5396_8177.n227 1.27228
R6807 a_5396_8177.n236 a_5396_8177.n233 1.27228
R6808 a_5396_8177.n188 a_5396_8177.n185 1.27228
R6809 a_5396_8177.n195 a_5396_8177.n192 1.27228
R6810 a_5396_8177.n201 a_5396_8177.n198 1.27228
R6811 a_5396_8177.n220 a_5396_8177.n214 1.27228
R6812 a_5396_8177.n176 a_5396_8177.n174 1.27228
R6813 a_5396_8177.n51 a_5396_8177.n50 1.26756
R6814 a_5396_8177.n63 a_5396_8177.n60 1.26756
R6815 a_5396_8177.n44 a_5396_8177.n43 1.26756
R6816 a_5396_8177.n275 a_5396_8177.n274 1.26756
R6817 a_5396_8177.n239 a_5396_8177.n238 1.15732
R6818 a_5396_8177.n205 a_5396_8177.n126 0.822966
R6819 a_5396_8177.n203 a_5396_8177.n202 0.822966
R6820 a_5396_8177.n70 a_5396_8177.n53 0.796291
R6821 a_5396_8177.n59 a_5396_8177.n57 0.796291
R6822 a_5396_8177.n265 a_5396_8177.n46 0.796291
R6823 a_5396_8177.n281 a_5396_8177.n277 0.796291
R6824 a_5396_8177.n100 a_5396_8177.n91 0.780703
R6825 a_5396_8177.n263 a_5396_8177.n242 0.780703
R6826 a_5396_8177.n283 a_5396_8177.n38 0.780703
R6827 a_5396_8177.n239 a_5396_8177.n39 0.780703
R6828 a_5396_8177.n223 a_5396_8177.n222 0.639318
R6829 a_5396_8177.n167 a_5396_8177.n126 0.639318
R6830 a_5396_8177.n237 a_5396_8177.n114 0.639318
R6831 a_5396_8177.n202 a_5396_8177.n177 0.639318
R6832 a_5396_8177.n264 a_5396_8177.n263 0.638405
R6833 a_5396_8177.n282 a_5396_8177.n39 0.638405
R6834 a_5396_8177.n264 a_5396_8177.n100 0.628372
R6835 a_5396_8177.n283 a_5396_8177.n282 0.628372
R6836 a_5396_8177.n222 a_5396_8177.n205 0.585196
R6837 a_5396_8177.n203 a_5396_8177.n114 0.585196
R6838 a_5396_8177.n70 a_5396_8177.n69 0.476484
R6839 a_5396_8177.n57 a_5396_8177.n56 0.476484
R6840 a_5396_8177.n268 a_5396_8177.n265 0.476484
R6841 a_5396_8177.n281 a_5396_8177.n280 0.476484
R6842 a_5396_8177.n241 a_5396_8177.n15 0.478684
R6843 a_5396_8177.n240 a_5396_8177.n9 0.478684
R6844 a_5396_8177.n99 a_5396_8177.n5 0.478684
R6845 a_5396_8177.n284 a_5396_8177.n0 0.478684
R6846 a_5396_8177.n224 a_5396_8177.n125 0.236091
R6847 a_5396_8177.n189 a_5396_8177.n188 0.236091
R6848 a_5396_8177.n17 a_5396_8177.n18 1.27228
R6849 a_5396_8177.n16 a_5396_8177.n17 2.51878
R6850 a_5396_8177.n241 a_5396_8177.n16 0.794091
R6851 a_5396_8177.n14 a_5396_8177.n15 1.27228
R6852 a_5396_8177.n13 a_5396_8177.n14 2.60203
R6853 a_5396_8177.n12 a_5396_8177.n13 1.27228
R6854 a_5396_8177.n11 a_5396_8177.n12 1.27228
R6855 a_5396_8177.n10 a_5396_8177.n11 2.51878
R6856 a_5396_8177.n240 a_5396_8177.n10 0.794091
R6857 a_5396_8177.t77 a_5396_8177.n9 6.77266
R6858 a_5396_8177.n24 a_5396_8177.n25 3.79678
R6859 a_5396_8177.n23 a_5396_8177.n24 1.27228
R6860 a_5396_8177.n204 a_5396_8177.n23 0.238291
R6861 a_5396_8177.n21 a_5396_8177.n22 1.27228
R6862 a_5396_8177.n20 a_5396_8177.n21 3.79678
R6863 a_5396_8177.n19 a_5396_8177.n20 1.27228
R6864 a_5396_8177.n203 a_5396_8177.n19 1.73829
R6865 a_5396_8177.n31 a_5396_8177.n32 3.79678
R6866 a_5396_8177.n30 a_5396_8177.n31 1.27228
R6867 a_5396_8177.n166 a_5396_8177.n30 0.238291
R6868 a_5396_8177.n28 a_5396_8177.n29 1.27228
R6869 a_5396_8177.n27 a_5396_8177.n28 3.79678
R6870 a_5396_8177.n26 a_5396_8177.n27 1.27228
R6871 a_5396_8177.n26 a_5396_8177.n177 2.32299
R6872 a_5396_8177.n7 a_5396_8177.n8 1.27228
R6873 a_5396_8177.n6 a_5396_8177.n7 2.51878
R6874 a_5396_8177.n99 a_5396_8177.n6 0.794091
R6875 a_5396_8177.n4 a_5396_8177.n5 1.27228
R6876 a_5396_8177.n3 a_5396_8177.n4 2.60203
R6877 a_5396_8177.n33 a_5396_8177.n3 1.27263
R6878 a_5396_8177.n33 a_5396_8177.n2 1.27192
R6879 a_5396_8177.n1 a_5396_8177.n2 2.51878
R6880 a_5396_8177.n284 a_5396_8177.n1 0.794091
R6881 a_5396_8177.t53 a_5396_8177.n0 6.77266
R6882 IREF.n1393 IREF.n1302 16.7377
R6883 IREF.n1303 IREF.t22 10.214
R6884 IREF.n1313 IREF.t50 10.214
R6885 IREF.n1324 IREF.t186 10.214
R6886 IREF.n1335 IREF.t110 10.214
R6887 IREF.n1346 IREF.t188 10.214
R6888 IREF.n1309 IREF.t8 10.2117
R6889 IREF.n1319 IREF.t147 10.2117
R6890 IREF.n1330 IREF.t55 10.2117
R6891 IREF.n1341 IREF.t210 10.2117
R6892 IREF.n1352 IREF.t57 10.2117
R6893 IREF.n1306 IREF.t218 9.58832
R6894 IREF.n1316 IREF.t123 9.58832
R6895 IREF.n1327 IREF.t2 9.58832
R6896 IREF.n1374 IREF.t243 9.58832
R6897 IREF.n1338 IREF.t16 9.58832
R6898 IREF.n1349 IREF.t260 9.58832
R6899 IREF.n1308 IREF.t259 9.58085
R6900 IREF.n1318 IREF.t175 9.58085
R6901 IREF.n1329 IREF.t34 9.58085
R6902 IREF.n1376 IREF.t69 9.58085
R6903 IREF.n1340 IREF.t6 9.58085
R6904 IREF.n1351 IREF.t91 9.58085
R6905 IREF.n1307 IREF.t250 9.58045
R6906 IREF.n1305 IREF.t28 9.58045
R6907 IREF.n1304 IREF.t40 9.58045
R6908 IREF.n1317 IREF.t165 9.58045
R6909 IREF.n1315 IREF.t242 9.58045
R6910 IREF.n1314 IREF.t208 9.58045
R6911 IREF.n1328 IREF.t38 9.58045
R6912 IREF.n1326 IREF.t151 9.58045
R6913 IREF.n1325 IREF.t111 9.58045
R6914 IREF.n1375 IREF.t54 9.58045
R6915 IREF.n1339 IREF.t12 9.58045
R6916 IREF.n1337 IREF.t83 9.58045
R6917 IREF.n1336 IREF.t263 9.58045
R6918 IREF.n1350 IREF.t82 9.58045
R6919 IREF.n1348 IREF.t155 9.58045
R6920 IREF.n1347 IREF.t112 9.58045
R6921 IREF.n1303 IREF.t42 9.58005
R6922 IREF.n1313 IREF.t194 9.58005
R6923 IREF.n1324 IREF.t101 9.58005
R6924 IREF.n1335 IREF.t252 9.58005
R6925 IREF.n1346 IREF.t104 9.58005
R6926 IREF.n1309 IREF.t32 9.57886
R6927 IREF.n1310 IREF.t20 9.57886
R6928 IREF.n1311 IREF.t10 9.57886
R6929 IREF.n1319 IREF.t237 9.57886
R6930 IREF.n1320 IREF.t77 9.57886
R6931 IREF.n1321 IREF.t135 9.57886
R6932 IREF.n1330 IREF.t139 9.57886
R6933 IREF.n1331 IREF.t209 9.57886
R6934 IREF.n1332 IREF.t271 9.57886
R6935 IREF.n1341 IREF.t67 9.57886
R6936 IREF.n1342 IREF.t126 9.57886
R6937 IREF.n1343 IREF.t199 9.57886
R6938 IREF.n1352 IREF.t140 9.57886
R6939 IREF.n1353 IREF.t212 9.57886
R6940 IREF.n1354 IREF.t44 9.57886
R6941 IREF.n1380 IREF.t0 8.38951
R6942 IREF.n1361 IREF.t18 8.38752
R6943 IREF.n833 IREF.t183 8.38704
R6944 IREF.n815 IREF.t166 8.38704
R6945 IREF.n947 IREF.t46 8.37857
R6946 IREF.n1070 IREF.t180 8.37857
R6947 IREF.n880 IREF.t214 8.31301
R6948 IREF.n1031 IREF.t115 8.31301
R6949 IREF.n1180 IREF.t264 8.29322
R6950 IREF.n969 IREF.t246 8.29322
R6951 IREF.n90 IREF.t255 8.10567
R6952 IREF.n1223 IREF.t244 8.10567
R6953 IREF.n1217 IREF.t95 8.10567
R6954 IREF.n1212 IREF.t192 8.10567
R6955 IREF.n1208 IREF.t207 8.10567
R6956 IREF.n1200 IREF.t117 8.10567
R6957 IREF.n134 IREF.t51 8.10567
R6958 IREF.n1270 IREF.t236 8.10567
R6959 IREF.n1276 IREF.t168 8.10567
R6960 IREF.n123 IREF.t160 8.10567
R6961 IREF.n116 IREF.t172 8.10567
R6962 IREF.n111 IREF.t45 8.10567
R6963 IREF.n1297 IREF.t58 8.10567
R6964 IREF.n1206 IREF.t62 8.10567
R6965 IREF.n1205 IREF.t227 8.10567
R6966 IREF.n1255 IREF.t70 8.10567
R6967 IREF.n104 IREF.t205 8.10567
R6968 IREF.n97 IREF.t132 8.10567
R6969 IREF.n55 IREF.t149 8.10567
R6970 IREF.n62 IREF.t176 8.10567
R6971 IREF.n64 IREF.t163 8.10567
R6972 IREF.n68 IREF.t145 8.10567
R6973 IREF.n219 IREF.t162 8.10567
R6974 IREF.n292 IREF.t72 8.10567
R6975 IREF.n286 IREF.t60 8.10567
R6976 IREF.n281 IREF.t215 8.10567
R6977 IREF.n276 IREF.t257 8.10567
R6978 IREF.n336 IREF.t105 8.10567
R6979 IREF.n346 IREF.t181 8.10567
R6980 IREF.n355 IREF.t86 8.10567
R6981 IREF.n364 IREF.t157 8.10567
R6982 IREF.n253 IREF.t225 8.10567
R6983 IREF.n246 IREF.t269 8.10567
R6984 IREF.n241 IREF.t198 8.10567
R6985 IREF.n236 IREF.t245 8.10567
R6986 IREF.n273 IREF.t64 8.10567
R6987 IREF.n272 IREF.t138 8.10567
R6988 IREF.n332 IREF.t127 8.10567
R6989 IREF.n233 IREF.t222 8.10567
R6990 IREF.n226 IREF.t68 8.10567
R6991 IREF.n176 IREF.t114 8.10567
R6992 IREF.n208 IREF.t167 8.10567
R6993 IREF.n199 IREF.t99 8.10567
R6994 IREF.n190 IREF.t234 8.10567
R6995 IREF.n406 IREF.t152 8.10567
R6996 IREF.n541 IREF.t53 8.10567
R6997 IREF.n535 IREF.t273 8.10567
R6998 IREF.n530 IREF.t202 8.10567
R6999 IREF.n559 IREF.t248 8.10567
R7000 IREF.n509 IREF.t96 8.10567
R7001 IREF.n153 IREF.t170 8.10567
R7002 IREF.n155 IREF.t74 8.10567
R7003 IREF.n486 IREF.t142 8.10567
R7004 IREF.n481 IREF.t211 8.10567
R7005 IREF.n165 IREF.t254 8.10567
R7006 IREF.n167 IREF.t182 8.10567
R7007 IREF.n458 IREF.t235 8.10567
R7008 IREF.n523 IREF.t258 8.10567
R7009 IREF.n516 IREF.t109 8.10567
R7010 IREF.n146 IREF.t103 8.10567
R7011 IREF.n454 IREF.t189 8.10567
R7012 IREF.n447 IREF.t262 8.10567
R7013 IREF.n404 IREF.t92 8.10567
R7014 IREF.n410 IREF.t156 8.10567
R7015 IREF.n415 IREF.t88 8.10567
R7016 IREF.n417 IREF.t221 8.10567
R7017 IREF.n601 IREF.t75 8.10567
R7018 IREF.n764 IREF.t203 8.10567
R7019 IREF.n758 IREF.t193 8.10567
R7020 IREF.n753 IREF.t119 8.10567
R7021 IREF.n748 IREF.t169 8.10567
R7022 IREF.n731 IREF.t240 8.10567
R7023 IREF.n720 IREF.t94 8.10567
R7024 IREF.n711 IREF.t219 8.10567
R7025 IREF.n702 IREF.t63 8.10567
R7026 IREF.n586 IREF.t124 8.10567
R7027 IREF.n682 IREF.t178 8.10567
R7028 IREF.n594 IREF.t102 8.10567
R7029 IREF.n598 IREF.t154 8.10567
R7030 IREF.n745 IREF.t197 8.10567
R7031 IREF.n738 IREF.t270 8.10567
R7032 IREF.n570 IREF.t261 8.10567
R7033 IREF.n647 IREF.t122 8.10567
R7034 IREF.n646 IREF.t201 8.10567
R7035 IREF.n657 IREF.t247 8.10567
R7036 IREF.n629 IREF.t80 8.10567
R7037 IREF.n609 IREF.t233 8.10567
R7038 IREF.n613 IREF.t131 8.10567
R7039 IREF.n1171 IREF.t134 8.10567
R7040 IREF.n1165 IREF.t78 8.10567
R7041 IREF.n1158 IREF.t251 8.10567
R7042 IREF.n802 IREF.t187 8.10567
R7043 IREF.n1175 IREF.t267 8.10567
R7044 IREF.n1174 IREF.t206 8.10567
R7045 IREF.n1173 IREF.t272 8.10567
R7046 IREF.n1179 IREF.t107 8.10567
R7047 IREF.n1185 IREF.t216 8.10567
R7048 IREF.n1191 IREF.t228 8.10567
R7049 IREF.n810 IREF.t49 8.10567
R7050 IREF.n812 IREF.t196 8.10567
R7051 IREF.n814 IREF.t185 8.10567
R7052 IREF.n1133 IREF.t184 8.10567
R7053 IREF.n1132 IREF.t116 8.10567
R7054 IREF.n1131 IREF.t125 8.10567
R7055 IREF.n1152 IREF.t179 8.10567
R7056 IREF.n1145 IREF.t190 8.10567
R7057 IREF.n806 IREF.t71 8.10567
R7058 IREF.n808 IREF.t85 8.10567
R7059 IREF.n938 IREF.t93 8.10567
R7060 IREF.n931 IREF.t161 8.10567
R7061 IREF.n925 IREF.t61 8.10567
R7062 IREF.n919 IREF.t133 8.10567
R7063 IREF.n942 IREF.t89 8.10567
R7064 IREF.n941 IREF.t159 8.10567
R7065 IREF.n940 IREF.t153 8.10567
R7066 IREF.n946 IREF.t265 8.10567
R7067 IREF.n945 IREF.t191 8.10567
R7068 IREF.n957 IREF.t241 8.10567
R7069 IREF.n875 IREF.t143 8.10567
R7070 IREF.n884 IREF.t146 8.10567
R7071 IREF.n879 IREF.t84 8.10567
R7072 IREF.n897 IREF.t238 8.10567
R7073 IREF.n896 IREF.t90 8.10567
R7074 IREF.n895 IREF.t130 8.10567
R7075 IREF.n917 IREF.t204 8.10567
R7076 IREF.n910 IREF.t249 8.10567
R7077 IREF.n903 IREF.t177 8.10567
R7078 IREF.n874 IREF.t232 8.10567
R7079 IREF.n861 IREF.t59 8.10567
R7080 IREF.n859 IREF.t129 8.10567
R7081 IREF.n858 IREF.t256 8.10567
R7082 IREF.n1002 IREF.t108 8.10567
R7083 IREF.n983 IREF.t76 8.10567
R7084 IREF.n984 IREF.t144 8.10567
R7085 IREF.n985 IREF.t136 8.10567
R7086 IREF.n968 IREF.t239 8.10567
R7087 IREF.n966 IREF.t164 8.10567
R7088 IREF.n965 IREF.t217 8.10567
R7089 IREF.n844 IREF.t113 8.10567
R7090 IREF.n838 IREF.t118 8.10567
R7091 IREF.n832 IREF.t47 8.10567
R7092 IREF.n848 IREF.t230 8.10567
R7093 IREF.n847 IREF.t81 8.10567
R7094 IREF.n846 IREF.t120 8.10567
R7095 IREF.n854 IREF.t174 8.10567
R7096 IREF.n853 IREF.t226 8.10567
R7097 IREF.n1014 IREF.t150 8.10567
R7098 IREF.n1020 IREF.t200 8.10567
R7099 IREF.n1064 IREF.t224 8.10567
R7100 IREF.n1060 IREF.t73 8.10567
R7101 IREF.n1059 IREF.t195 8.10567
R7102 IREF.n1103 IREF.t268 8.10567
R7103 IREF.n1083 IREF.t220 8.10567
R7104 IREF.n1084 IREF.t65 8.10567
R7105 IREF.n1085 IREF.t56 8.10567
R7106 IREF.n1069 IREF.t173 8.10567
R7107 IREF.n1067 IREF.t100 8.10567
R7108 IREF.n1065 IREF.t148 8.10567
R7109 IREF.n1045 IREF.t48 8.10567
R7110 IREF.n1038 IREF.t52 8.10567
R7111 IREF.n1032 IREF.t213 8.10567
R7112 IREF.n1049 IREF.t141 8.10567
R7113 IREF.n1048 IREF.t223 8.10567
R7114 IREF.n1047 IREF.t266 8.10567
R7115 IREF.n1105 IREF.t106 8.10567
R7116 IREF.n1053 IREF.t158 8.10567
R7117 IREF.n1052 IREF.t87 8.10567
R7118 IREF.n1122 IREF.t128 8.10567
R7119 IREF.n1381 IREF.t26 8.10567
R7120 IREF.n1386 IREF.t14 8.10567
R7121 IREF.n1377 IREF.t4 8.10567
R7122 IREF.n1372 IREF.t24 8.10567
R7123 IREF.n1365 IREF.t30 8.10567
R7124 IREF.n1360 IREF.t36 8.10567
R7125 IREF.n27 IREF.n24 6.61324
R7126 IREF.n35 IREF.t9 6.47665
R7127 IREF.n7 IREF.n6 6.43481
R7128 IREF.n23 IREF.t1 6.43476
R7129 IREF.n30 IREF.n29 5.34147
R7130 IREF.n28 IREF.t29 5.34147
R7131 IREF.n192 IREF.n189 4.65575
R7132 IREF.n614 IREF.n612 4.65575
R7133 IREF.n293 IREF.n290 4.64641
R7134 IREF.n765 IREF.n760 4.64641
R7135 IREF.n1153 IREF.n1152 4.64261
R7136 IREF.n1004 IREF.n854 4.64261
R7137 IREF.n1373 IREF.n1372 4.64261
R7138 IREF.n69 IREF.n67 4.64
R7139 IREF.n1225 IREF.n1224 4.64
R7140 IREF.n296 IREF.n290 4.64
R7141 IREF.n418 IREF.n416 4.64
R7142 IREF.n543 IREF.n542 4.64
R7143 IREF.n420 IREF.n416 4.64
R7144 IREF.n544 IREF.n543 4.64
R7145 IREF.n766 IREF.n765 4.64
R7146 IREF.n70 IREF.n69 4.64
R7147 IREF.n1226 IREF.n1225 4.64
R7148 IREF.n918 IREF.n917 4.61892
R7149 IREF.n1106 IREF.n1105 4.61892
R7150 IREF.n920 IREF.n919 4.61655
R7151 IREF.n1104 IREF.n1103 4.61655
R7152 IREF.n35 IREF.n34 4.61078
R7153 IREF.n21 IREF.n20 4.61078
R7154 IREF.n16 IREF.n15 4.61078
R7155 IREF.n12 IREF.n11 4.61078
R7156 IREF.n23 IREF.n2 4.61078
R7157 IREF.n45 IREF.n43 4.60951
R7158 IREF.n46 IREF.n45 4.60951
R7159 IREF.n20 IREF.n17 4.60825
R7160 IREF.n15 IREF.n13 4.60825
R7161 IREF.n11 IREF.n7 4.60825
R7162 IREF.n22 IREF.n2 4.60825
R7163 IREF.n1245 IREF.n1206 4.54125
R7164 IREF.n105 IREF.n104 4.54125
R7165 IREF.n524 IREF.n523 4.54125
R7166 IREF.n455 IREF.n454 4.54125
R7167 IREF.n322 IREF.n273 4.53893
R7168 IREF.n234 IREF.n233 4.53893
R7169 IREF.n746 IREF.n745 4.53893
R7170 IREF.n647 IREF.n599 4.53893
R7171 IREF.n320 IREF.n275 4.51011
R7172 IREF.n367 IREF.n366 4.51011
R7173 IREF.n397 IREF.n396 4.51011
R7174 IREF.n792 IREF.n791 4.51011
R7175 IREF.n699 IREF.n584 4.51011
R7176 IREF.n665 IREF.n663 4.51011
R7177 IREF.n335 IREF.n267 4.50691
R7178 IREF.n369 IREF.n368 4.50691
R7179 IREF.n220 IREF.n170 4.50691
R7180 IREF.n732 IREF.n564 4.50691
R7181 IREF.n698 IREF.n697 4.50691
R7182 IREF.n661 IREF.n660 4.50691
R7183 IREF.n44 IREF.n37 4.5005
R7184 IREF.n103 IREF.n52 4.5005
R7185 IREF.n102 IREF.n101 4.5005
R7186 IREF.n100 IREF.n53 4.5005
R7187 IREF.n99 IREF.n98 4.5005
R7188 IREF.n96 IREF.n54 4.5005
R7189 IREF.n95 IREF.n94 4.5005
R7190 IREF.n1247 IREF.n1246 4.5005
R7191 IREF.n1248 IREF.n1204 4.5005
R7192 IREF.n1250 IREF.n1249 4.5005
R7193 IREF.n1251 IREF.n1203 4.5005
R7194 IREF.n1253 IREF.n1252 4.5005
R7195 IREF.n1254 IREF.n1202 4.5005
R7196 IREF.n1280 IREF.n1279 4.5005
R7197 IREF.n124 IREF.n121 4.5005
R7198 IREF.n1284 IREF.n120 4.5005
R7199 IREF.n1285 IREF.n119 4.5005
R7200 IREF.n1286 IREF.n118 4.5005
R7201 IREF.n1289 IREF.n115 4.5005
R7202 IREF.n1290 IREF.n114 4.5005
R7203 IREF.n1291 IREF.n113 4.5005
R7204 IREF.n112 IREF.n109 4.5005
R7205 IREF.n1295 IREF.n108 4.5005
R7206 IREF.n1296 IREF.n107 4.5005
R7207 IREF.n1298 IREF.n106 4.5005
R7208 IREF.n1258 IREF.n1257 4.5005
R7209 IREF.n1201 IREF.n139 4.5005
R7210 IREF.n1262 IREF.n138 4.5005
R7211 IREF.n1263 IREF.n137 4.5005
R7212 IREF.n1264 IREF.n136 4.5005
R7213 IREF.n135 IREF.n132 4.5005
R7214 IREF.n1268 IREF.n131 4.5005
R7215 IREF.n1269 IREF.n130 4.5005
R7216 IREF.n1271 IREF.n129 4.5005
R7217 IREF.n128 IREF.n126 4.5005
R7218 IREF.n1275 IREF.n125 4.5005
R7219 IREF.n1278 IREF.n1277 4.5005
R7220 IREF.n1224 IREF.n1222 4.5005
R7221 IREF.n1228 IREF.n1221 4.5005
R7222 IREF.n1229 IREF.n1220 4.5005
R7223 IREF.n1230 IREF.n1219 4.5005
R7224 IREF.n1233 IREF.n1216 4.5005
R7225 IREF.n1234 IREF.n1215 4.5005
R7226 IREF.n1235 IREF.n1214 4.5005
R7227 IREF.n1238 IREF.n1211 4.5005
R7228 IREF.n1239 IREF.n1210 4.5005
R7229 IREF.n1240 IREF.n1207 4.5005
R7230 IREF.n1244 IREF.n1243 4.5005
R7231 IREF.n92 IREF.n91 4.5005
R7232 IREF.n89 IREF.n56 4.5005
R7233 IREF.n83 IREF.n57 4.5005
R7234 IREF.n85 IREF.n84 4.5005
R7235 IREF.n82 IREF.n59 4.5005
R7236 IREF.n81 IREF.n80 4.5005
R7237 IREF.n61 IREF.n60 4.5005
R7238 IREF.n76 IREF.n75 4.5005
R7239 IREF.n74 IREF.n73 4.5005
R7240 IREF.n72 IREF.n65 4.5005
R7241 IREF.n67 IREF.n66 4.5005
R7242 IREF.n232 IREF.n173 4.5005
R7243 IREF.n231 IREF.n230 4.5005
R7244 IREF.n229 IREF.n174 4.5005
R7245 IREF.n228 IREF.n227 4.5005
R7246 IREF.n225 IREF.n175 4.5005
R7247 IREF.n224 IREF.n223 4.5005
R7248 IREF.n324 IREF.n323 4.5005
R7249 IREF.n325 IREF.n271 4.5005
R7250 IREF.n327 IREF.n326 4.5005
R7251 IREF.n328 IREF.n270 4.5005
R7252 IREF.n330 IREF.n329 4.5005
R7253 IREF.n331 IREF.n269 4.5005
R7254 IREF.n396 IREF.n395 4.5005
R7255 IREF.n394 IREF.n393 4.5005
R7256 IREF.n237 IREF.n235 4.5005
R7257 IREF.n388 IREF.n387 4.5005
R7258 IREF.n386 IREF.n385 4.5005
R7259 IREF.n242 IREF.n240 4.5005
R7260 IREF.n380 IREF.n379 4.5005
R7261 IREF.n378 IREF.n377 4.5005
R7262 IREF.n247 IREF.n245 4.5005
R7263 IREF.n251 IREF.n249 4.5005
R7264 IREF.n372 IREF.n371 4.5005
R7265 IREF.n370 IREF.n369 4.5005
R7266 IREF.n366 IREF.n252 4.5005
R7267 IREF.n363 IREF.n362 4.5005
R7268 IREF.n361 IREF.n360 4.5005
R7269 IREF.n257 IREF.n256 4.5005
R7270 IREF.n354 IREF.n353 4.5005
R7271 IREF.n352 IREF.n351 4.5005
R7272 IREF.n262 IREF.n261 4.5005
R7273 IREF.n345 IREF.n344 4.5005
R7274 IREF.n343 IREF.n342 4.5005
R7275 IREF.n341 IREF.n265 4.5005
R7276 IREF.n268 IREF.n266 4.5005
R7277 IREF.n335 IREF.n334 4.5005
R7278 IREF.n321 IREF.n320 4.5005
R7279 IREF.n278 IREF.n274 4.5005
R7280 IREF.n315 IREF.n314 4.5005
R7281 IREF.n313 IREF.n312 4.5005
R7282 IREF.n283 IREF.n280 4.5005
R7283 IREF.n307 IREF.n306 4.5005
R7284 IREF.n305 IREF.n304 4.5005
R7285 IREF.n288 IREF.n285 4.5005
R7286 IREF.n299 IREF.n298 4.5005
R7287 IREF.n297 IREF.n289 4.5005
R7288 IREF.n296 IREF.n295 4.5005
R7289 IREF.n192 IREF.n191 4.5005
R7290 IREF.n194 IREF.n193 4.5005
R7291 IREF.n186 IREF.n185 4.5005
R7292 IREF.n201 IREF.n200 4.5005
R7293 IREF.n203 IREF.n202 4.5005
R7294 IREF.n182 IREF.n181 4.5005
R7295 IREF.n211 IREF.n210 4.5005
R7296 IREF.n212 IREF.n180 4.5005
R7297 IREF.n214 IREF.n213 4.5005
R7298 IREF.n178 IREF.n177 4.5005
R7299 IREF.n221 IREF.n220 4.5005
R7300 IREF.n188 IREF.n187 4.5005
R7301 IREF.n196 IREF.n195 4.5005
R7302 IREF.n198 IREF.n197 4.5005
R7303 IREF.n184 IREF.n183 4.5005
R7304 IREF.n205 IREF.n204 4.5005
R7305 IREF.n207 IREF.n206 4.5005
R7306 IREF.n209 IREF.n179 4.5005
R7307 IREF.n216 IREF.n215 4.5005
R7308 IREF.n218 IREF.n217 4.5005
R7309 IREF.n172 IREF.n171 4.5005
R7310 IREF.n392 IREF.n391 4.5005
R7311 IREF.n390 IREF.n389 4.5005
R7312 IREF.n239 IREF.n238 4.5005
R7313 IREF.n384 IREF.n383 4.5005
R7314 IREF.n382 IREF.n381 4.5005
R7315 IREF.n244 IREF.n243 4.5005
R7316 IREF.n376 IREF.n375 4.5005
R7317 IREF.n374 IREF.n373 4.5005
R7318 IREF.n250 IREF.n248 4.5005
R7319 IREF.n365 IREF.n254 4.5005
R7320 IREF.n258 IREF.n255 4.5005
R7321 IREF.n359 IREF.n358 4.5005
R7322 IREF.n357 IREF.n356 4.5005
R7323 IREF.n260 IREF.n259 4.5005
R7324 IREF.n350 IREF.n349 4.5005
R7325 IREF.n348 IREF.n347 4.5005
R7326 IREF.n264 IREF.n263 4.5005
R7327 IREF.n340 IREF.n339 4.5005
R7328 IREF.n338 IREF.n337 4.5005
R7329 IREF.n319 IREF.n318 4.5005
R7330 IREF.n317 IREF.n316 4.5005
R7331 IREF.n279 IREF.n277 4.5005
R7332 IREF.n311 IREF.n310 4.5005
R7333 IREF.n309 IREF.n308 4.5005
R7334 IREF.n284 IREF.n282 4.5005
R7335 IREF.n303 IREF.n302 4.5005
R7336 IREF.n301 IREF.n300 4.5005
R7337 IREF.n291 IREF.n287 4.5005
R7338 IREF.n294 IREF.n293 4.5005
R7339 IREF.n453 IREF.n401 4.5005
R7340 IREF.n452 IREF.n451 4.5005
R7341 IREF.n450 IREF.n402 4.5005
R7342 IREF.n449 IREF.n448 4.5005
R7343 IREF.n446 IREF.n403 4.5005
R7344 IREF.n445 IREF.n444 4.5005
R7345 IREF.n522 IREF.n143 4.5005
R7346 IREF.n521 IREF.n520 4.5005
R7347 IREF.n519 IREF.n144 4.5005
R7348 IREF.n518 IREF.n517 4.5005
R7349 IREF.n515 IREF.n145 4.5005
R7350 IREF.n514 IREF.n513 4.5005
R7351 IREF.n483 IREF.n482 4.5005
R7352 IREF.n480 IREF.n159 4.5005
R7353 IREF.n474 IREF.n160 4.5005
R7354 IREF.n476 IREF.n475 4.5005
R7355 IREF.n473 IREF.n162 4.5005
R7356 IREF.n472 IREF.n471 4.5005
R7357 IREF.n164 IREF.n163 4.5005
R7358 IREF.n467 IREF.n466 4.5005
R7359 IREF.n465 IREF.n464 4.5005
R7360 IREF.n463 IREF.n168 4.5005
R7361 IREF.n456 IREF.n169 4.5005
R7362 IREF.n459 IREF.n457 4.5005
R7363 IREF.n511 IREF.n510 4.5005
R7364 IREF.n508 IREF.n147 4.5005
R7365 IREF.n502 IREF.n148 4.5005
R7366 IREF.n504 IREF.n503 4.5005
R7367 IREF.n501 IREF.n150 4.5005
R7368 IREF.n500 IREF.n499 4.5005
R7369 IREF.n152 IREF.n151 4.5005
R7370 IREF.n495 IREF.n494 4.5005
R7371 IREF.n493 IREF.n492 4.5005
R7372 IREF.n491 IREF.n156 4.5005
R7373 IREF.n484 IREF.n157 4.5005
R7374 IREF.n487 IREF.n485 4.5005
R7375 IREF.n542 IREF.n540 4.5005
R7376 IREF.n546 IREF.n539 4.5005
R7377 IREF.n547 IREF.n538 4.5005
R7378 IREF.n548 IREF.n537 4.5005
R7379 IREF.n551 IREF.n534 4.5005
R7380 IREF.n552 IREF.n533 4.5005
R7381 IREF.n553 IREF.n532 4.5005
R7382 IREF.n531 IREF.n528 4.5005
R7383 IREF.n557 IREF.n527 4.5005
R7384 IREF.n558 IREF.n526 4.5005
R7385 IREF.n560 IREF.n525 4.5005
R7386 IREF.n442 IREF.n441 4.5005
R7387 IREF.n438 IREF.n405 4.5005
R7388 IREF.n437 IREF.n436 4.5005
R7389 IREF.n435 IREF.n408 4.5005
R7390 IREF.n434 IREF.n433 4.5005
R7391 IREF.n429 IREF.n409 4.5005
R7392 IREF.n428 IREF.n427 4.5005
R7393 IREF.n426 IREF.n412 4.5005
R7394 IREF.n425 IREF.n424 4.5005
R7395 IREF.n414 IREF.n413 4.5005
R7396 IREF.n419 IREF.n418 4.5005
R7397 IREF.n420 IREF.n419 4.5005
R7398 IREF.n421 IREF.n414 4.5005
R7399 IREF.n424 IREF.n423 4.5005
R7400 IREF.n422 IREF.n412 4.5005
R7401 IREF.n428 IREF.n411 4.5005
R7402 IREF.n430 IREF.n429 4.5005
R7403 IREF.n433 IREF.n432 4.5005
R7404 IREF.n431 IREF.n408 4.5005
R7405 IREF.n437 IREF.n407 4.5005
R7406 IREF.n439 IREF.n438 4.5005
R7407 IREF.n441 IREF.n440 4.5005
R7408 IREF.n460 IREF.n459 4.5005
R7409 IREF.n461 IREF.n169 4.5005
R7410 IREF.n463 IREF.n462 4.5005
R7411 IREF.n464 IREF.n166 4.5005
R7412 IREF.n468 IREF.n467 4.5005
R7413 IREF.n469 IREF.n164 4.5005
R7414 IREF.n471 IREF.n470 4.5005
R7415 IREF.n162 IREF.n161 4.5005
R7416 IREF.n477 IREF.n476 4.5005
R7417 IREF.n478 IREF.n160 4.5005
R7418 IREF.n480 IREF.n479 4.5005
R7419 IREF.n482 IREF.n158 4.5005
R7420 IREF.n488 IREF.n487 4.5005
R7421 IREF.n489 IREF.n157 4.5005
R7422 IREF.n491 IREF.n490 4.5005
R7423 IREF.n492 IREF.n154 4.5005
R7424 IREF.n496 IREF.n495 4.5005
R7425 IREF.n497 IREF.n152 4.5005
R7426 IREF.n499 IREF.n498 4.5005
R7427 IREF.n150 IREF.n149 4.5005
R7428 IREF.n505 IREF.n504 4.5005
R7429 IREF.n506 IREF.n148 4.5005
R7430 IREF.n508 IREF.n507 4.5005
R7431 IREF.n510 IREF.n141 4.5005
R7432 IREF.n561 IREF.n560 4.5005
R7433 IREF.n558 IREF.n142 4.5005
R7434 IREF.n557 IREF.n556 4.5005
R7435 IREF.n555 IREF.n528 4.5005
R7436 IREF.n554 IREF.n553 4.5005
R7437 IREF.n552 IREF.n529 4.5005
R7438 IREF.n551 IREF.n550 4.5005
R7439 IREF.n549 IREF.n548 4.5005
R7440 IREF.n547 IREF.n536 4.5005
R7441 IREF.n546 IREF.n545 4.5005
R7442 IREF.n544 IREF.n540 4.5005
R7443 IREF.n649 IREF.n648 4.5005
R7444 IREF.n650 IREF.n645 4.5005
R7445 IREF.n652 IREF.n651 4.5005
R7446 IREF.n653 IREF.n644 4.5005
R7447 IREF.n655 IREF.n654 4.5005
R7448 IREF.n656 IREF.n643 4.5005
R7449 IREF.n744 IREF.n567 4.5005
R7450 IREF.n743 IREF.n742 4.5005
R7451 IREF.n741 IREF.n568 4.5005
R7452 IREF.n740 IREF.n739 4.5005
R7453 IREF.n737 IREF.n569 4.5005
R7454 IREF.n736 IREF.n735 4.5005
R7455 IREF.n666 IREF.n665 4.5005
R7456 IREF.n668 IREF.n667 4.5005
R7457 IREF.n596 IREF.n595 4.5005
R7458 IREF.n675 IREF.n674 4.5005
R7459 IREF.n677 IREF.n676 4.5005
R7460 IREF.n592 IREF.n591 4.5005
R7461 IREF.n685 IREF.n684 4.5005
R7462 IREF.n686 IREF.n590 4.5005
R7463 IREF.n688 IREF.n687 4.5005
R7464 IREF.n588 IREF.n587 4.5005
R7465 IREF.n695 IREF.n694 4.5005
R7466 IREF.n697 IREF.n696 4.5005
R7467 IREF.n584 IREF.n583 4.5005
R7468 IREF.n704 IREF.n703 4.5005
R7469 IREF.n706 IREF.n705 4.5005
R7470 IREF.n580 IREF.n579 4.5005
R7471 IREF.n713 IREF.n712 4.5005
R7472 IREF.n715 IREF.n714 4.5005
R7473 IREF.n576 IREF.n575 4.5005
R7474 IREF.n723 IREF.n722 4.5005
R7475 IREF.n724 IREF.n574 4.5005
R7476 IREF.n726 IREF.n725 4.5005
R7477 IREF.n572 IREF.n571 4.5005
R7478 IREF.n733 IREF.n732 4.5005
R7479 IREF.n791 IREF.n790 4.5005
R7480 IREF.n789 IREF.n788 4.5005
R7481 IREF.n749 IREF.n747 4.5005
R7482 IREF.n783 IREF.n782 4.5005
R7483 IREF.n781 IREF.n780 4.5005
R7484 IREF.n754 IREF.n752 4.5005
R7485 IREF.n775 IREF.n774 4.5005
R7486 IREF.n773 IREF.n772 4.5005
R7487 IREF.n759 IREF.n757 4.5005
R7488 IREF.n763 IREF.n761 4.5005
R7489 IREF.n767 IREF.n766 4.5005
R7490 IREF.n615 IREF.n614 4.5005
R7491 IREF.n611 IREF.n610 4.5005
R7492 IREF.n622 IREF.n621 4.5005
R7493 IREF.n624 IREF.n623 4.5005
R7494 IREF.n607 IREF.n606 4.5005
R7495 IREF.n632 IREF.n631 4.5005
R7496 IREF.n633 IREF.n605 4.5005
R7497 IREF.n635 IREF.n634 4.5005
R7498 IREF.n603 IREF.n602 4.5005
R7499 IREF.n642 IREF.n641 4.5005
R7500 IREF.n660 IREF.n659 4.5005
R7501 IREF.n617 IREF.n616 4.5005
R7502 IREF.n619 IREF.n618 4.5005
R7503 IREF.n620 IREF.n608 4.5005
R7504 IREF.n626 IREF.n625 4.5005
R7505 IREF.n628 IREF.n627 4.5005
R7506 IREF.n630 IREF.n604 4.5005
R7507 IREF.n637 IREF.n636 4.5005
R7508 IREF.n639 IREF.n638 4.5005
R7509 IREF.n640 IREF.n600 4.5005
R7510 IREF.n664 IREF.n597 4.5005
R7511 IREF.n670 IREF.n669 4.5005
R7512 IREF.n672 IREF.n671 4.5005
R7513 IREF.n673 IREF.n593 4.5005
R7514 IREF.n679 IREF.n678 4.5005
R7515 IREF.n681 IREF.n680 4.5005
R7516 IREF.n683 IREF.n589 4.5005
R7517 IREF.n690 IREF.n689 4.5005
R7518 IREF.n692 IREF.n691 4.5005
R7519 IREF.n693 IREF.n585 4.5005
R7520 IREF.n701 IREF.n700 4.5005
R7521 IREF.n582 IREF.n581 4.5005
R7522 IREF.n708 IREF.n707 4.5005
R7523 IREF.n710 IREF.n709 4.5005
R7524 IREF.n578 IREF.n577 4.5005
R7525 IREF.n717 IREF.n716 4.5005
R7526 IREF.n719 IREF.n718 4.5005
R7527 IREF.n721 IREF.n573 4.5005
R7528 IREF.n728 IREF.n727 4.5005
R7529 IREF.n730 IREF.n729 4.5005
R7530 IREF.n566 IREF.n565 4.5005
R7531 IREF.n787 IREF.n786 4.5005
R7532 IREF.n785 IREF.n784 4.5005
R7533 IREF.n751 IREF.n750 4.5005
R7534 IREF.n779 IREF.n778 4.5005
R7535 IREF.n777 IREF.n776 4.5005
R7536 IREF.n756 IREF.n755 4.5005
R7537 IREF.n771 IREF.n770 4.5005
R7538 IREF.n769 IREF.n768 4.5005
R7539 IREF.n762 IREF.n760 4.5005
R7540 IREF.n70 IREF.n66 4.5005
R7541 IREF.n72 IREF.n71 4.5005
R7542 IREF.n73 IREF.n63 4.5005
R7543 IREF.n77 IREF.n76 4.5005
R7544 IREF.n78 IREF.n61 4.5005
R7545 IREF.n80 IREF.n79 4.5005
R7546 IREF.n59 IREF.n58 4.5005
R7547 IREF.n86 IREF.n85 4.5005
R7548 IREF.n87 IREF.n57 4.5005
R7549 IREF.n89 IREF.n88 4.5005
R7550 IREF.n91 IREF.n50 4.5005
R7551 IREF.n1299 IREF.n1298 4.5005
R7552 IREF.n1296 IREF.n51 4.5005
R7553 IREF.n1295 IREF.n1294 4.5005
R7554 IREF.n1293 IREF.n109 4.5005
R7555 IREF.n1292 IREF.n1291 4.5005
R7556 IREF.n1290 IREF.n110 4.5005
R7557 IREF.n1289 IREF.n1288 4.5005
R7558 IREF.n1287 IREF.n1286 4.5005
R7559 IREF.n1285 IREF.n117 4.5005
R7560 IREF.n1284 IREF.n1283 4.5005
R7561 IREF.n1282 IREF.n121 4.5005
R7562 IREF.n1281 IREF.n1280 4.5005
R7563 IREF.n1277 IREF.n122 4.5005
R7564 IREF.n1275 IREF.n1274 4.5005
R7565 IREF.n1273 IREF.n126 4.5005
R7566 IREF.n1272 IREF.n1271 4.5005
R7567 IREF.n1269 IREF.n127 4.5005
R7568 IREF.n1268 IREF.n1267 4.5005
R7569 IREF.n1266 IREF.n132 4.5005
R7570 IREF.n1265 IREF.n1264 4.5005
R7571 IREF.n1263 IREF.n133 4.5005
R7572 IREF.n1262 IREF.n1261 4.5005
R7573 IREF.n1260 IREF.n139 4.5005
R7574 IREF.n1259 IREF.n1258 4.5005
R7575 IREF.n1243 IREF.n1242 4.5005
R7576 IREF.n1241 IREF.n1240 4.5005
R7577 IREF.n1239 IREF.n1209 4.5005
R7578 IREF.n1238 IREF.n1237 4.5005
R7579 IREF.n1236 IREF.n1235 4.5005
R7580 IREF.n1234 IREF.n1213 4.5005
R7581 IREF.n1233 IREF.n1232 4.5005
R7582 IREF.n1231 IREF.n1230 4.5005
R7583 IREF.n1229 IREF.n1218 4.5005
R7584 IREF.n1228 IREF.n1227 4.5005
R7585 IREF.n1226 IREF.n1222 4.5005
R7586 IREF.n882 IREF.n881 4.5005
R7587 IREF.n883 IREF.n878 4.5005
R7588 IREF.n886 IREF.n885 4.5005
R7589 IREF.n887 IREF.n877 4.5005
R7590 IREF.n889 IREF.n888 4.5005
R7591 IREF.n890 IREF.n876 4.5005
R7592 IREF.n892 IREF.n891 4.5005
R7593 IREF.n894 IREF.n893 4.5005
R7594 IREF.n899 IREF.n898 4.5005
R7595 IREF.n901 IREF.n900 4.5005
R7596 IREF.n902 IREF.n873 4.5005
R7597 IREF.n905 IREF.n904 4.5005
R7598 IREF.n906 IREF.n872 4.5005
R7599 IREF.n908 IREF.n907 4.5005
R7600 IREF.n909 IREF.n871 4.5005
R7601 IREF.n912 IREF.n911 4.5005
R7602 IREF.n913 IREF.n870 4.5005
R7603 IREF.n915 IREF.n914 4.5005
R7604 IREF.n916 IREF.n869 4.5005
R7605 IREF.n921 IREF.n868 4.5005
R7606 IREF.n923 IREF.n922 4.5005
R7607 IREF.n924 IREF.n867 4.5005
R7608 IREF.n927 IREF.n926 4.5005
R7609 IREF.n928 IREF.n866 4.5005
R7610 IREF.n930 IREF.n929 4.5005
R7611 IREF.n932 IREF.n865 4.5005
R7612 IREF.n934 IREF.n933 4.5005
R7613 IREF.n935 IREF.n864 4.5005
R7614 IREF.n937 IREF.n936 4.5005
R7615 IREF.n939 IREF.n862 4.5005
R7616 IREF.n959 IREF.n958 4.5005
R7617 IREF.n956 IREF.n863 4.5005
R7618 IREF.n955 IREF.n954 4.5005
R7619 IREF.n953 IREF.n943 4.5005
R7620 IREF.n952 IREF.n951 4.5005
R7621 IREF.n950 IREF.n944 4.5005
R7622 IREF.n949 IREF.n948 4.5005
R7623 IREF.n845 IREF.n827 4.5005
R7624 IREF.n843 IREF.n842 4.5005
R7625 IREF.n841 IREF.n829 4.5005
R7626 IREF.n840 IREF.n839 4.5005
R7627 IREF.n837 IREF.n830 4.5005
R7628 IREF.n836 IREF.n835 4.5005
R7629 IREF.n834 IREF.n831 4.5005
R7630 IREF.n1023 IREF.n1022 4.5005
R7631 IREF.n1021 IREF.n828 4.5005
R7632 IREF.n1019 IREF.n1018 4.5005
R7633 IREF.n1017 IREF.n849 4.5005
R7634 IREF.n1016 IREF.n1015 4.5005
R7635 IREF.n1013 IREF.n850 4.5005
R7636 IREF.n1012 IREF.n1011 4.5005
R7637 IREF.n1010 IREF.n851 4.5005
R7638 IREF.n1009 IREF.n1008 4.5005
R7639 IREF.n1007 IREF.n852 4.5005
R7640 IREF.n1006 IREF.n1005 4.5005
R7641 IREF.n987 IREF.n986 4.5005
R7642 IREF.n989 IREF.n988 4.5005
R7643 IREF.n990 IREF.n860 4.5005
R7644 IREF.n992 IREF.n991 4.5005
R7645 IREF.n994 IREF.n993 4.5005
R7646 IREF.n995 IREF.n857 4.5005
R7647 IREF.n997 IREF.n996 4.5005
R7648 IREF.n998 IREF.n856 4.5005
R7649 IREF.n1000 IREF.n999 4.5005
R7650 IREF.n1001 IREF.n855 4.5005
R7651 IREF.n982 IREF.n981 4.5005
R7652 IREF.n980 IREF.n963 4.5005
R7653 IREF.n979 IREF.n978 4.5005
R7654 IREF.n977 IREF.n964 4.5005
R7655 IREF.n976 IREF.n975 4.5005
R7656 IREF.n974 IREF.n973 4.5005
R7657 IREF.n972 IREF.n967 4.5005
R7658 IREF.n971 IREF.n970 4.5005
R7659 IREF.n1034 IREF.n1033 4.5005
R7660 IREF.n1035 IREF.n1030 4.5005
R7661 IREF.n1037 IREF.n1036 4.5005
R7662 IREF.n1039 IREF.n1029 4.5005
R7663 IREF.n1041 IREF.n1040 4.5005
R7664 IREF.n1042 IREF.n1028 4.5005
R7665 IREF.n1044 IREF.n1043 4.5005
R7666 IREF.n1046 IREF.n1026 4.5005
R7667 IREF.n1124 IREF.n1123 4.5005
R7668 IREF.n1121 IREF.n1027 4.5005
R7669 IREF.n1120 IREF.n1119 4.5005
R7670 IREF.n1118 IREF.n1050 4.5005
R7671 IREF.n1117 IREF.n1116 4.5005
R7672 IREF.n1115 IREF.n1051 4.5005
R7673 IREF.n1114 IREF.n1113 4.5005
R7674 IREF.n1112 IREF.n1111 4.5005
R7675 IREF.n1110 IREF.n1054 4.5005
R7676 IREF.n1109 IREF.n1108 4.5005
R7677 IREF.n1107 IREF.n1055 4.5005
R7678 IREF.n1102 IREF.n1056 4.5005
R7679 IREF.n1101 IREF.n1100 4.5005
R7680 IREF.n1099 IREF.n1057 4.5005
R7681 IREF.n1098 IREF.n1097 4.5005
R7682 IREF.n1096 IREF.n1058 4.5005
R7683 IREF.n1095 IREF.n1094 4.5005
R7684 IREF.n1093 IREF.n1092 4.5005
R7685 IREF.n1091 IREF.n1061 4.5005
R7686 IREF.n1090 IREF.n1089 4.5005
R7687 IREF.n1088 IREF.n1062 4.5005
R7688 IREF.n1087 IREF.n1086 4.5005
R7689 IREF.n1082 IREF.n1081 4.5005
R7690 IREF.n1080 IREF.n1079 4.5005
R7691 IREF.n1078 IREF.n1066 4.5005
R7692 IREF.n1077 IREF.n1076 4.5005
R7693 IREF.n1075 IREF.n1074 4.5005
R7694 IREF.n1073 IREF.n1068 4.5005
R7695 IREF.n1072 IREF.n1071 4.5005
R7696 IREF.n1130 IREF.n1129 4.5005
R7697 IREF.n825 IREF.n824 4.5005
R7698 IREF.n823 IREF.n811 4.5005
R7699 IREF.n822 IREF.n821 4.5005
R7700 IREF.n820 IREF.n819 4.5005
R7701 IREF.n818 IREF.n813 4.5005
R7702 IREF.n817 IREF.n816 4.5005
R7703 IREF.n1134 IREF.n809 4.5005
R7704 IREF.n1136 IREF.n1135 4.5005
R7705 IREF.n1138 IREF.n1137 4.5005
R7706 IREF.n1139 IREF.n807 4.5005
R7707 IREF.n1141 IREF.n1140 4.5005
R7708 IREF.n1143 IREF.n1142 4.5005
R7709 IREF.n1144 IREF.n805 4.5005
R7710 IREF.n1147 IREF.n1146 4.5005
R7711 IREF.n1148 IREF.n804 4.5005
R7712 IREF.n1150 IREF.n1149 4.5005
R7713 IREF.n1151 IREF.n803 4.5005
R7714 IREF.n1172 IREF.n796 4.5005
R7715 IREF.n1170 IREF.n1169 4.5005
R7716 IREF.n1168 IREF.n798 4.5005
R7717 IREF.n1167 IREF.n1166 4.5005
R7718 IREF.n1164 IREF.n799 4.5005
R7719 IREF.n1163 IREF.n1162 4.5005
R7720 IREF.n1161 IREF.n800 4.5005
R7721 IREF.n1160 IREF.n1159 4.5005
R7722 IREF.n1157 IREF.n801 4.5005
R7723 IREF.n1156 IREF.n1155 4.5005
R7724 IREF.n1194 IREF.n1193 4.5005
R7725 IREF.n1192 IREF.n797 4.5005
R7726 IREF.n1190 IREF.n1189 4.5005
R7727 IREF.n1188 IREF.n1176 4.5005
R7728 IREF.n1187 IREF.n1186 4.5005
R7729 IREF.n1184 IREF.n1177 4.5005
R7730 IREF.n1183 IREF.n1182 4.5005
R7731 IREF.n1181 IREF.n1178 4.5005
R7732 IREF.n1363 IREF.n1362 4.5005
R7733 IREF.n1364 IREF.n1359 4.5005
R7734 IREF.n1367 IREF.n1366 4.5005
R7735 IREF.n1368 IREF.n1358 4.5005
R7736 IREF.n1370 IREF.n1369 4.5005
R7737 IREF.n1371 IREF.n1357 4.5005
R7738 IREF.n1389 IREF.n1388 4.5005
R7739 IREF.n1387 IREF.n1378 4.5005
R7740 IREF.n1386 IREF.n1385 4.5005
R7741 IREF.n1384 IREF.n1379 4.5005
R7742 IREF.n1383 IREF.n1382 4.5005
R7743 IREF.n10 IREF.n5 4.5005
R7744 IREF.n14 IREF.n4 4.5005
R7745 IREF.n19 IREF.n3 4.5005
R7746 IREF.n1397 IREF.n1396 4.5005
R7747 IREF.n1197 IREF.n48 3.97759
R7748 IREF.n27 IREF.n26 3.87147
R7749 IREF.n44 IREF.t35 3.86699
R7750 IREF.n19 IREF.n18 3.83383
R7751 IREF.n14 IREF.t25 3.83383
R7752 IREF.n45 IREF.t7 3.66094
R7753 IREF.n1004 IREF.n1003 3.03856
R7754 IREF.n1154 IREF.n1153 3.03856
R7755 IREF.n1279 IREF.n1278 3.0245
R7756 IREF.n370 IREF.n252 3.0245
R7757 IREF.n485 IREF.n483 3.0245
R7758 IREF.n488 IREF.n158 3.0245
R7759 IREF.n696 IREF.n583 3.0245
R7760 IREF.n1281 IREF.n122 3.0245
R7761 IREF.n920 IREF.n918 3.0245
R7762 IREF.n1106 IREF.n1104 3.0245
R7763 IREF.n368 IREF.n367 2.96825
R7764 IREF.n699 IREF.n698 2.96825
R7765 IREF.n47 IREF.n46 2.94838
R7766 IREF.n43 IREF.n42 2.60059
R7767 IREF.n30 IREF.n28 2.51878
R7768 IREF.n47 IREF.n36 2.44398
R7769 IREF.n189 IREF.n187 2.41967
R7770 IREF.n617 IREF.n612 2.41967
R7771 IREF.n34 IREF.n33 2.40646
R7772 IREF.n42 IREF.n39 2.39895
R7773 IREF.n10 IREF.n9 2.36383
R7774 IREF.n1025 IREF.n826 2.30989
R7775 IREF.n961 IREF.n960 2.30989
R7776 IREF IREF.n1 2.28212
R7777 IREF.n1154 IREF.n802 2.25752
R7778 IREF.n1003 IREF.n1002 2.25752
R7779 IREF.n1390 IREF.n1377 2.25278
R7780 IREF.n17 IREF.n16 2.246
R7781 IREF.n34 IREF.n31 2.24358
R7782 IREF.n1256 IREF.n1255 2.22849
R7783 IREF.n93 IREF.n55 2.22849
R7784 IREF.n512 IREF.n146 2.22849
R7785 IREF.n443 IREF.n404 2.22849
R7786 IREF.n333 IREF.n332 2.22782
R7787 IREF.n222 IREF.n176 2.22782
R7788 IREF.n734 IREF.n570 2.22782
R7789 IREF.n658 IREF.n657 2.22782
R7790 IREF.n42 IREF.n41 2.19216
R7791 IREF.n893 IREF.n826 2.18975
R7792 IREF.n960 IREF.n862 2.18975
R7793 IREF.n1125 IREF.n1026 2.18975
R7794 IREF.n1087 IREF.n1063 2.18975
R7795 IREF.n1024 IREF.n827 2.16725
R7796 IREF.n987 IREF.n962 2.16725
R7797 IREF.n1129 IREF.n1128 2.16725
R7798 IREF.n1195 IREF.n796 2.16725
R7799 IREF.n460 IREF.n400 2.102
R7800 IREF.n562 IREF.n561 2.102
R7801 IREF.n1300 IREF.n1299 2.102
R7802 IREF.n1242 IREF.n1199 2.102
R7803 IREF.n399 IREF.n398 2.07182
R7804 IREF.n563 IREF.n140 2.07182
R7805 IREF.n398 IREF.n397 2.06825
R7806 IREF.n275 IREF.n140 2.06825
R7807 IREF.n663 IREF.n662 2.06825
R7808 IREF.n793 IREF.n792 2.06825
R7809 IREF.n1197 IREF.n1196 2.01366
R7810 IREF.n1394 IREF.n1393 1.91821
R7811 IREF.n1323 IREF.n1312 1.61908
R7812 IREF.n1302 IREF.n1301 1.53101
R7813 IREF.n1198 IREF.n1197 1.53101
R7814 IREF.n662 IREF.n49 1.5005
R7815 IREF.n400 IREF.n399 1.5005
R7816 IREF.n1301 IREF.n1300 1.5005
R7817 IREF.n1199 IREF.n1198 1.5005
R7818 IREF.n794 IREF.n793 1.5005
R7819 IREF.n563 IREF.n562 1.5005
R7820 IREF.n1126 IREF.n1125 1.5005
R7821 IREF.n1025 IREF.n1024 1.5005
R7822 IREF.n1128 IREF.n1127 1.5005
R7823 IREF.n1196 IREF.n1195 1.5005
R7824 IREF.n1063 IREF.n795 1.5005
R7825 IREF.n962 IREF.n961 1.5005
R7826 IREF.n1356 IREF.n1355 1.5005
R7827 IREF.n1345 IREF.n1344 1.5005
R7828 IREF.n1392 IREF.n1391 1.5005
R7829 IREF.n1334 IREF.n1333 1.5005
R7830 IREF.n1323 IREF.n1322 1.5005
R7831 IREF.n1395 IREF.n1394 1.5005
R7832 IREF.n399 IREF.n49 1.47516
R7833 IREF.n794 IREF.n563 1.47516
R7834 IREF.n1 IREF.t15 1.4705
R7835 IREF.n1 IREF.n0 1.4705
R7836 IREF.n33 IREF.t21 1.4705
R7837 IREF.n33 IREF.n32 1.4705
R7838 IREF.n26 IREF.t43 1.4705
R7839 IREF.n26 IREF.n25 1.4705
R7840 IREF.n39 IREF.t3 1.4705
R7841 IREF.n39 IREF.n38 1.4705
R7842 IREF.n41 IREF.t17 1.4705
R7843 IREF.n41 IREF.n40 1.4705
R7844 IREF.n9 IREF.t37 1.4705
R7845 IREF.n9 IREF.n8 1.4705
R7846 IREF.n1393 IREF.n1392 1.42915
R7847 IREF.n1127 IREF.n48 1.41182
R7848 IREF.n970 IREF.n969 1.392
R7849 IREF.n1181 IREF.n1180 1.392
R7850 IREF.n881 IREF.n880 1.38741
R7851 IREF.n1034 IREF.n1031 1.38741
R7852 IREF.n28 IREF.n27 1.27228
R7853 IREF.n958 IREF.n942 1.24866
R7854 IREF.n898 IREF.n897 1.24866
R7855 IREF.n1083 IREF.n1082 1.24866
R7856 IREF.n1123 IREF.n1049 1.24866
R7857 IREF.n940 IREF.n939 1.24629
R7858 IREF.n895 IREF.n894 1.24629
R7859 IREF.n1086 IREF.n1085 1.24629
R7860 IREF.n1047 IREF.n1046 1.24629
R7861 IREF.n1126 IREF.n1025 1.23709
R7862 IREF.n961 IREF.n795 1.23709
R7863 IREF.n1173 IREF.n1172 1.22261
R7864 IREF.n1131 IREF.n1130 1.22261
R7865 IREF.n986 IREF.n985 1.22261
R7866 IREF.n846 IREF.n845 1.22261
R7867 IREF.n1193 IREF.n1175 1.21313
R7868 IREF.n1134 IREF.n1133 1.21313
R7869 IREF.n983 IREF.n982 1.21313
R7870 IREF.n1022 IREF.n848 1.21313
R7871 IREF.n31 IREF.n30 1.20609
R7872 IREF.n834 IREF.n833 1.12904
R7873 IREF.n816 IREF.n815 1.12904
R7874 IREF.n1362 IREF.n1361 1.129
R7875 IREF.n1383 IREF.n1380 1.12765
R7876 IREF.n948 IREF.n947 1.11862
R7877 IREF.n1071 IREF.n1070 1.11862
R7878 IREF.n13 IREF.n12 0.9995
R7879 IREF.n22 IREF.n21 0.9995
R7880 IREF.n1306 IREF.n1305 0.915282
R7881 IREF.n1316 IREF.n1315 0.915282
R7882 IREF.n1327 IREF.n1326 0.915282
R7883 IREF.n1338 IREF.n1337 0.915282
R7884 IREF.n1349 IREF.n1348 0.915282
R7885 IREF.n1394 IREF.n47 0.886209
R7886 IREF.n440 IREF.n400 0.83975
R7887 IREF.n562 IREF.n141 0.83975
R7888 IREF.n1300 IREF.n50 0.83975
R7889 IREF.n1259 IREF.n1199 0.83975
R7890 IREF.n398 IREF.n170 0.81725
R7891 IREF.n267 IREF.n140 0.81725
R7892 IREF.n662 IREF.n661 0.81725
R7893 IREF.n793 IREF.n564 0.81725
R7894 IREF.n1127 IREF.n1126 0.809892
R7895 IREF.n1196 IREF.n795 0.809892
R7896 IREF.n1374 IREF.n1373 0.779178
R7897 IREF.n93 IREF.n92 0.75626
R7898 IREF.n1257 IREF.n1256 0.75626
R7899 IREF.n443 IREF.n442 0.75626
R7900 IREF.n512 IREF.n511 0.75626
R7901 IREF.n222 IREF.n221 0.756242
R7902 IREF.n334 IREF.n333 0.756242
R7903 IREF.n659 IREF.n658 0.756242
R7904 IREF.n734 IREF.n733 0.756242
R7905 IREF.n899 IREF.n826 0.752
R7906 IREF.n960 IREF.n959 0.752
R7907 IREF.n1125 IREF.n1124 0.752
R7908 IREF.n1081 IREF.n1063 0.752
R7909 IREF.n1024 IREF.n1023 0.71825
R7910 IREF.n981 IREF.n962 0.71825
R7911 IREF.n1128 IREF.n809 0.71825
R7912 IREF.n1195 IREF.n1194 0.71825
R7913 IREF.n106 IREF.n105 0.698
R7914 IREF.n1245 IREF.n1244 0.698
R7915 IREF.n395 IREF.n234 0.698
R7916 IREF.n322 IREF.n321 0.698
R7917 IREF.n457 IREF.n455 0.698
R7918 IREF.n525 IREF.n524 0.698
R7919 IREF.n666 IREF.n599 0.698
R7920 IREF.n790 IREF.n746 0.698
R7921 IREF.n1312 IREF.n1311 0.688348
R7922 IREF.n1322 IREF.n1321 0.688348
R7923 IREF.n1333 IREF.n1332 0.688348
R7924 IREF.n1344 IREF.n1343 0.688348
R7925 IREF.n1355 IREF.n1354 0.688348
R7926 IREF.n1174 IREF.n1173 0.673132
R7927 IREF.n1175 IREF.n1174 0.673132
R7928 IREF.n1132 IREF.n1131 0.673132
R7929 IREF.n1133 IREF.n1132 0.673132
R7930 IREF.n941 IREF.n940 0.673132
R7931 IREF.n942 IREF.n941 0.673132
R7932 IREF.n896 IREF.n895 0.673132
R7933 IREF.n897 IREF.n896 0.673132
R7934 IREF.n985 IREF.n984 0.673132
R7935 IREF.n984 IREF.n983 0.673132
R7936 IREF.n847 IREF.n846 0.673132
R7937 IREF.n848 IREF.n847 0.673132
R7938 IREF.n1085 IREF.n1084 0.673132
R7939 IREF.n1084 IREF.n1083 0.673132
R7940 IREF.n1048 IREF.n1047 0.673132
R7941 IREF.n1049 IREF.n1048 0.673132
R7942 IREF.n1307 IREF.n1306 0.655148
R7943 IREF.n1317 IREF.n1316 0.655148
R7944 IREF.n1328 IREF.n1327 0.655148
R7945 IREF.n1375 IREF.n1374 0.655148
R7946 IREF.n1339 IREF.n1338 0.655148
R7947 IREF.n1350 IREF.n1349 0.655148
R7948 IREF.n1305 IREF.n1304 0.63334
R7949 IREF.n1311 IREF.n1310 0.63334
R7950 IREF.n1310 IREF.n1309 0.63334
R7951 IREF.n1315 IREF.n1314 0.63334
R7952 IREF.n1321 IREF.n1320 0.63334
R7953 IREF.n1320 IREF.n1319 0.63334
R7954 IREF.n1326 IREF.n1325 0.63334
R7955 IREF.n1332 IREF.n1331 0.63334
R7956 IREF.n1331 IREF.n1330 0.63334
R7957 IREF.n1337 IREF.n1336 0.63334
R7958 IREF.n1343 IREF.n1342 0.63334
R7959 IREF.n1342 IREF.n1341 0.63334
R7960 IREF.n1348 IREF.n1347 0.63334
R7961 IREF.n1354 IREF.n1353 0.63334
R7962 IREF.n1353 IREF.n1352 0.63334
R7963 IREF.n1304 IREF.n1303 0.63225
R7964 IREF.n1308 IREF.n1307 0.63225
R7965 IREF.n1314 IREF.n1313 0.63225
R7966 IREF.n1318 IREF.n1317 0.63225
R7967 IREF.n1325 IREF.n1324 0.63225
R7968 IREF.n1329 IREF.n1328 0.63225
R7969 IREF.n1376 IREF.n1375 0.63225
R7970 IREF.n1336 IREF.n1335 0.63225
R7971 IREF.n1340 IREF.n1339 0.63225
R7972 IREF.n1347 IREF.n1346 0.63225
R7973 IREF.n1351 IREF.n1350 0.63225
R7974 IREF.n1391 IREF.n1390 0.622055
R7975 IREF.n1302 IREF.n48 0.602344
R7976 IREF.n1301 IREF.n49 0.571818
R7977 IREF.n1198 IREF.n794 0.571818
R7978 IREF.n1345 IREF.n1334 0.467527
R7979 IREF.n1180 IREF.n1179 0.45279
R7980 IREF.n969 IREF.n968 0.45279
R7981 IREF.n880 IREF.n879 0.430924
R7982 IREF.n1032 IREF.n1031 0.430924
R7983 IREF.n950 IREF.n949 0.394842
R7984 IREF.n930 IREF.n866 0.394842
R7985 IREF.n909 IREF.n908 0.394842
R7986 IREF.n885 IREF.n883 0.394842
R7987 IREF.n1073 IREF.n1072 0.394842
R7988 IREF.n1096 IREF.n1095 0.394842
R7989 IREF.n1115 IREF.n1114 0.394842
R7990 IREF.n1037 IREF.n1030 0.394842
R7991 IREF.n955 IREF.n943 0.381816
R7992 IREF.n924 IREF.n923 0.381816
R7993 IREF.n904 IREF.n902 0.381816
R7994 IREF.n1078 IREF.n1077 0.381816
R7995 IREF.n1101 IREF.n1057 0.381816
R7996 IREF.n1120 IREF.n1050 0.381816
R7997 IREF.n1190 IREF.n1176 0.379447
R7998 IREF.n1184 IREF.n1183 0.379447
R7999 IREF.n1157 IREF.n1156 0.379447
R8000 IREF.n1163 IREF.n800 0.379447
R8001 IREF.n1166 IREF.n798 0.379447
R8002 IREF.n1139 IREF.n1138 0.379447
R8003 IREF.n1144 IREF.n1143 0.379447
R8004 IREF.n1150 IREF.n804 0.379447
R8005 IREF.n818 IREF.n817 0.379447
R8006 IREF.n823 IREF.n822 0.379447
R8007 IREF.n978 IREF.n977 0.379447
R8008 IREF.n973 IREF.n972 0.379447
R8009 IREF.n1001 IREF.n1000 0.379447
R8010 IREF.n996 IREF.n995 0.379447
R8011 IREF.n991 IREF.n990 0.379447
R8012 IREF.n1019 IREF.n849 0.379447
R8013 IREF.n1013 IREF.n1012 0.379447
R8014 IREF.n1008 IREF.n1007 0.379447
R8015 IREF.n836 IREF.n831 0.379447
R8016 IREF.n839 IREF.n829 0.379447
R8017 IREF.n1388 IREF.n1387 0.379447
R8018 IREF.n1382 IREF.n1379 0.379447
R8019 IREF.n1370 IREF.n1358 0.379447
R8020 IREF.n1364 IREF.n1363 0.378263
R8021 IREF.n81 IREF.n60 0.375125
R8022 IREF.n115 IREF.n114 0.375125
R8023 IREF.n135 IREF.n131 0.375125
R8024 IREF.n1216 IREF.n1215 0.375125
R8025 IREF.n202 IREF.n181 0.375125
R8026 IREF.n379 IREF.n240 0.375125
R8027 IREF.n352 IREF.n261 0.375125
R8028 IREF.n306 IREF.n305 0.375125
R8029 IREF.n427 IREF.n409 0.375125
R8030 IREF.n472 IREF.n163 0.375125
R8031 IREF.n500 IREF.n151 0.375125
R8032 IREF.n534 IREF.n533 0.375125
R8033 IREF.n430 IREF.n411 0.375125
R8034 IREF.n470 IREF.n469 0.375125
R8035 IREF.n498 IREF.n497 0.375125
R8036 IREF.n550 IREF.n529 0.375125
R8037 IREF.n632 IREF.n606 0.375125
R8038 IREF.n685 IREF.n591 0.375125
R8039 IREF.n714 IREF.n575 0.375125
R8040 IREF.n774 IREF.n752 0.375125
R8041 IREF.n79 IREF.n78 0.375125
R8042 IREF.n1288 IREF.n110 0.375125
R8043 IREF.n1267 IREF.n1266 0.375125
R8044 IREF.n1232 IREF.n1213 0.375125
R8045 IREF.n886 IREF.n878 0.375125
R8046 IREF.n907 IREF.n871 0.375125
R8047 IREF.n929 IREF.n928 0.375125
R8048 IREF.n948 IREF.n944 0.375125
R8049 IREF.n1036 IREF.n1035 0.375125
R8050 IREF.n1113 IREF.n1051 0.375125
R8051 IREF.n1094 IREF.n1058 0.375125
R8052 IREF.n1071 IREF.n1068 0.375125
R8053 IREF.n74 IREF.n65 0.36275
R8054 IREF.n112 IREF.n108 0.36275
R8055 IREF.n129 IREF.n128 0.36275
R8056 IREF.n1211 IREF.n1210 0.36275
R8057 IREF.n193 IREF.n185 0.36275
R8058 IREF.n387 IREF.n235 0.36275
R8059 IREF.n361 IREF.n256 0.36275
R8060 IREF.n314 IREF.n313 0.36275
R8061 IREF.n425 IREF.n413 0.36275
R8062 IREF.n465 IREF.n168 0.36275
R8063 IREF.n493 IREF.n156 0.36275
R8064 IREF.n531 IREF.n527 0.36275
R8065 IREF.n423 IREF.n421 0.36275
R8066 IREF.n462 IREF.n166 0.36275
R8067 IREF.n490 IREF.n154 0.36275
R8068 IREF.n556 IREF.n555 0.36275
R8069 IREF.n622 IREF.n610 0.36275
R8070 IREF.n675 IREF.n595 0.36275
R8071 IREF.n705 IREF.n579 0.36275
R8072 IREF.n782 IREF.n747 0.36275
R8073 IREF.n71 IREF.n63 0.36275
R8074 IREF.n1294 IREF.n1293 0.36275
R8075 IREF.n1273 IREF.n1272 0.36275
R8076 IREF.n1237 IREF.n1209 0.36275
R8077 IREF.n905 IREF.n873 0.36275
R8078 IREF.n922 IREF.n867 0.36275
R8079 IREF.n954 IREF.n953 0.36275
R8080 IREF.n1119 IREF.n1118 0.36275
R8081 IREF.n1100 IREF.n1099 0.36275
R8082 IREF.n1076 IREF.n1066 0.36275
R8083 IREF.n94 IREF.n54 0.3605
R8084 IREF.n101 IREF.n100 0.3605
R8085 IREF.n1252 IREF.n1202 0.3605
R8086 IREF.n1250 IREF.n1204 0.3605
R8087 IREF.n223 IREF.n175 0.3605
R8088 IREF.n230 IREF.n229 0.3605
R8089 IREF.n329 IREF.n269 0.3605
R8090 IREF.n327 IREF.n271 0.3605
R8091 IREF.n196 IREF.n187 0.3605
R8092 IREF.n205 IREF.n183 0.3605
R8093 IREF.n216 IREF.n179 0.3605
R8094 IREF.n391 IREF.n390 0.3605
R8095 IREF.n383 IREF.n382 0.3605
R8096 IREF.n375 IREF.n374 0.3605
R8097 IREF.n358 IREF.n258 0.3605
R8098 IREF.n349 IREF.n259 0.3605
R8099 IREF.n339 IREF.n263 0.3605
R8100 IREF.n317 IREF.n277 0.3605
R8101 IREF.n309 IREF.n282 0.3605
R8102 IREF.n301 IREF.n287 0.3605
R8103 IREF.n444 IREF.n403 0.3605
R8104 IREF.n451 IREF.n450 0.3605
R8105 IREF.n513 IREF.n145 0.3605
R8106 IREF.n520 IREF.n519 0.3605
R8107 IREF.n654 IREF.n643 0.3605
R8108 IREF.n652 IREF.n645 0.3605
R8109 IREF.n735 IREF.n569 0.3605
R8110 IREF.n742 IREF.n741 0.3605
R8111 IREF.n618 IREF.n617 0.3605
R8112 IREF.n627 IREF.n626 0.3605
R8113 IREF.n638 IREF.n637 0.3605
R8114 IREF.n671 IREF.n670 0.3605
R8115 IREF.n680 IREF.n679 0.3605
R8116 IREF.n691 IREF.n690 0.3605
R8117 IREF.n708 IREF.n581 0.3605
R8118 IREF.n717 IREF.n577 0.3605
R8119 IREF.n728 IREF.n573 0.3605
R8120 IREF.n786 IREF.n785 0.3605
R8121 IREF.n778 IREF.n777 0.3605
R8122 IREF.n770 IREF.n769 0.3605
R8123 IREF.n835 IREF.n834 0.3605
R8124 IREF.n841 IREF.n840 0.3605
R8125 IREF.n1018 IREF.n1017 0.3605
R8126 IREF.n1011 IREF.n850 0.3605
R8127 IREF.n1009 IREF.n852 0.3605
R8128 IREF.n999 IREF.n855 0.3605
R8129 IREF.n997 IREF.n857 0.3605
R8130 IREF.n992 IREF.n860 0.3605
R8131 IREF.n979 IREF.n964 0.3605
R8132 IREF.n974 IREF.n967 0.3605
R8133 IREF.n816 IREF.n813 0.3605
R8134 IREF.n821 IREF.n811 0.3605
R8135 IREF.n1137 IREF.n807 0.3605
R8136 IREF.n1142 IREF.n805 0.3605
R8137 IREF.n1149 IREF.n1148 0.3605
R8138 IREF.n1155 IREF.n801 0.3605
R8139 IREF.n1162 IREF.n1161 0.3605
R8140 IREF.n1168 IREF.n1167 0.3605
R8141 IREF.n1189 IREF.n1188 0.3605
R8142 IREF.n1182 IREF.n1177 0.3605
R8143 IREF.n1369 IREF.n1368 0.3605
R8144 IREF.n1389 IREF.n1378 0.3605
R8145 IREF.n1384 IREF.n1383 0.3605
R8146 IREF.n1362 IREF.n1359 0.359375
R8147 IREF.n947 IREF.n946 0.348488
R8148 IREF.n1070 IREF.n1069 0.348488
R8149 IREF.n815 IREF.n814 0.327481
R8150 IREF.n833 IREF.n832 0.327481
R8151 IREF.n1361 IREF.n1360 0.32675
R8152 IREF.n1381 IREF.n1380 0.324133
R8153 IREF.n1356 IREF.n1345 0.307291
R8154 IREF.n933 IREF.n864 0.302474
R8155 IREF.n915 IREF.n870 0.302474
R8156 IREF.n890 IREF.n889 0.302474
R8157 IREF.n1091 IREF.n1090 0.302474
R8158 IREF.n1110 IREF.n1109 0.302474
R8159 IREF.n1040 IREF.n1028 0.302474
R8160 IREF.n1334 IREF.n1323 0.301209
R8161 IREF.n84 IREF.n83 0.287375
R8162 IREF.n120 IREF.n119 0.287375
R8163 IREF.n138 IREF.n137 0.287375
R8164 IREF.n1221 IREF.n1220 0.287375
R8165 IREF.n213 IREF.n212 0.287375
R8166 IREF.n251 IREF.n245 0.287375
R8167 IREF.n343 IREF.n265 0.287375
R8168 IREF.n298 IREF.n297 0.287375
R8169 IREF.n436 IREF.n435 0.287375
R8170 IREF.n475 IREF.n474 0.287375
R8171 IREF.n503 IREF.n502 0.287375
R8172 IREF.n539 IREF.n538 0.287375
R8173 IREF.n431 IREF.n407 0.287375
R8174 IREF.n478 IREF.n477 0.287375
R8175 IREF.n506 IREF.n505 0.287375
R8176 IREF.n545 IREF.n536 0.287375
R8177 IREF.n634 IREF.n602 0.287375
R8178 IREF.n687 IREF.n587 0.287375
R8179 IREF.n725 IREF.n724 0.287375
R8180 IREF.n763 IREF.n757 0.287375
R8181 IREF.n87 IREF.n86 0.287375
R8182 IREF.n1283 IREF.n117 0.287375
R8183 IREF.n1261 IREF.n133 0.287375
R8184 IREF.n1227 IREF.n1218 0.287375
R8185 IREF.n888 IREF.n876 0.287375
R8186 IREF.n914 IREF.n913 0.287375
R8187 IREF.n935 IREF.n934 0.287375
R8188 IREF.n1042 IREF.n1041 0.287375
R8189 IREF.n1108 IREF.n1054 0.287375
R8190 IREF.n1089 IREF.n1061 0.287375
R8191 IREF.n1312 IREF.n1308 0.254694
R8192 IREF.n1322 IREF.n1318 0.254694
R8193 IREF.n1333 IREF.n1329 0.254694
R8194 IREF.n1391 IREF.n1376 0.254694
R8195 IREF.n1344 IREF.n1340 0.254694
R8196 IREF.n1355 IREF.n1351 0.254694
R8197 IREF.n223 IREF.n222 0.208888
R8198 IREF.n333 IREF.n269 0.208888
R8199 IREF.n658 IREF.n643 0.208888
R8200 IREF.n735 IREF.n734 0.208888
R8201 IREF.n94 IREF.n93 0.20887
R8202 IREF.n1256 IREF.n1202 0.20887
R8203 IREF.n444 IREF.n443 0.20887
R8204 IREF.n513 IREF.n512 0.20887
R8205 IREF.n1003 IREF.n855 0.208099
R8206 IREF.n1155 IREF.n1154 0.208099
R8207 IREF.n1390 IREF.n1389 0.208099
R8208 IREF.n1193 IREF.n1192 0.147342
R8209 IREF.n1186 IREF.n1176 0.147342
R8210 IREF.n1183 IREF.n1178 0.147342
R8211 IREF.n1159 IREF.n1157 0.147342
R8212 IREF.n1164 IREF.n1163 0.147342
R8213 IREF.n1170 IREF.n798 0.147342
R8214 IREF.n1135 IREF.n1134 0.147342
R8215 IREF.n1140 IREF.n1139 0.147342
R8216 IREF.n1146 IREF.n1144 0.147342
R8217 IREF.n1151 IREF.n1150 0.147342
R8218 IREF.n819 IREF.n818 0.147342
R8219 IREF.n824 IREF.n823 0.147342
R8220 IREF.n956 IREF.n955 0.147342
R8221 IREF.n951 IREF.n950 0.147342
R8222 IREF.n923 IREF.n868 0.147342
R8223 IREF.n926 IREF.n866 0.147342
R8224 IREF.n933 IREF.n932 0.147342
R8225 IREF.n937 IREF.n864 0.147342
R8226 IREF.n902 IREF.n901 0.147342
R8227 IREF.n908 IREF.n872 0.147342
R8228 IREF.n911 IREF.n870 0.147342
R8229 IREF.n916 IREF.n915 0.147342
R8230 IREF.n883 IREF.n882 0.147342
R8231 IREF.n889 IREF.n877 0.147342
R8232 IREF.n891 IREF.n890 0.147342
R8233 IREF.n982 IREF.n963 0.147342
R8234 IREF.n977 IREF.n976 0.147342
R8235 IREF.n972 IREF.n971 0.147342
R8236 IREF.n1000 IREF.n856 0.147342
R8237 IREF.n995 IREF.n994 0.147342
R8238 IREF.n990 IREF.n989 0.147342
R8239 IREF.n1022 IREF.n1021 0.147342
R8240 IREF.n1015 IREF.n849 0.147342
R8241 IREF.n1012 IREF.n851 0.147342
R8242 IREF.n1007 IREF.n1006 0.147342
R8243 IREF.n837 IREF.n836 0.147342
R8244 IREF.n843 IREF.n829 0.147342
R8245 IREF.n1079 IREF.n1078 0.147342
R8246 IREF.n1074 IREF.n1073 0.147342
R8247 IREF.n1102 IREF.n1101 0.147342
R8248 IREF.n1097 IREF.n1096 0.147342
R8249 IREF.n1092 IREF.n1091 0.147342
R8250 IREF.n1090 IREF.n1062 0.147342
R8251 IREF.n1121 IREF.n1120 0.147342
R8252 IREF.n1116 IREF.n1115 0.147342
R8253 IREF.n1111 IREF.n1110 0.147342
R8254 IREF.n1109 IREF.n1055 0.147342
R8255 IREF.n1033 IREF.n1030 0.147342
R8256 IREF.n1040 IREF.n1039 0.147342
R8257 IREF.n1044 IREF.n1028 0.147342
R8258 IREF.n1388 IREF.n1377 0.147342
R8259 IREF.n1387 IREF.n1386 0.147342
R8260 IREF.n1386 IREF.n1379 0.147342
R8261 IREF.n1382 IREF.n1381 0.147342
R8262 IREF.n1366 IREF.n1364 0.147342
R8263 IREF.n1371 IREF.n1370 0.147342
R8264 IREF.n1363 IREF.n1360 0.143789
R8265 IREF.n1191 IREF.n1190 0.142605
R8266 IREF.n1185 IREF.n1184 0.142605
R8267 IREF.n1156 IREF.n802 0.142605
R8268 IREF.n1158 IREF.n800 0.142605
R8269 IREF.n1166 IREF.n1165 0.142605
R8270 IREF.n1172 IREF.n1171 0.142605
R8271 IREF.n1138 IREF.n808 0.142605
R8272 IREF.n1143 IREF.n806 0.142605
R8273 IREF.n1145 IREF.n804 0.142605
R8274 IREF.n817 IREF.n814 0.142605
R8275 IREF.n822 IREF.n812 0.142605
R8276 IREF.n1130 IREF.n810 0.142605
R8277 IREF.n978 IREF.n965 0.142605
R8278 IREF.n973 IREF.n966 0.142605
R8279 IREF.n1002 IREF.n1001 0.142605
R8280 IREF.n996 IREF.n858 0.142605
R8281 IREF.n991 IREF.n859 0.142605
R8282 IREF.n986 IREF.n861 0.142605
R8283 IREF.n1020 IREF.n1019 0.142605
R8284 IREF.n1014 IREF.n1013 0.142605
R8285 IREF.n1008 IREF.n853 0.142605
R8286 IREF.n832 IREF.n831 0.142605
R8287 IREF.n839 IREF.n838 0.142605
R8288 IREF.n845 IREF.n844 0.142605
R8289 IREF.n1365 IREF.n1358 0.142605
R8290 IREF.n43 IREF.n37 0.14
R8291 IREF.n46 IREF.n37 0.14
R8292 IREF.n67 IREF.n65 0.14
R8293 IREF.n75 IREF.n74 0.14
R8294 IREF.n75 IREF.n60 0.14
R8295 IREF.n82 IREF.n81 0.14
R8296 IREF.n84 IREF.n82 0.14
R8297 IREF.n83 IREF.n56 0.14
R8298 IREF.n92 IREF.n56 0.14
R8299 IREF.n99 IREF.n54 0.14
R8300 IREF.n100 IREF.n99 0.14
R8301 IREF.n101 IREF.n52 0.14
R8302 IREF.n105 IREF.n52 0.14
R8303 IREF.n107 IREF.n106 0.14
R8304 IREF.n108 IREF.n107 0.14
R8305 IREF.n113 IREF.n112 0.14
R8306 IREF.n114 IREF.n113 0.14
R8307 IREF.n118 IREF.n115 0.14
R8308 IREF.n119 IREF.n118 0.14
R8309 IREF.n124 IREF.n120 0.14
R8310 IREF.n1279 IREF.n124 0.14
R8311 IREF.n1278 IREF.n125 0.14
R8312 IREF.n128 IREF.n125 0.14
R8313 IREF.n130 IREF.n129 0.14
R8314 IREF.n131 IREF.n130 0.14
R8315 IREF.n136 IREF.n135 0.14
R8316 IREF.n137 IREF.n136 0.14
R8317 IREF.n1201 IREF.n138 0.14
R8318 IREF.n1257 IREF.n1201 0.14
R8319 IREF.n1252 IREF.n1251 0.14
R8320 IREF.n1251 IREF.n1250 0.14
R8321 IREF.n1246 IREF.n1204 0.14
R8322 IREF.n1246 IREF.n1245 0.14
R8323 IREF.n1244 IREF.n1207 0.14
R8324 IREF.n1210 IREF.n1207 0.14
R8325 IREF.n1214 IREF.n1211 0.14
R8326 IREF.n1215 IREF.n1214 0.14
R8327 IREF.n1219 IREF.n1216 0.14
R8328 IREF.n1220 IREF.n1219 0.14
R8329 IREF.n1224 IREF.n1221 0.14
R8330 IREF.n193 IREF.n192 0.14
R8331 IREF.n201 IREF.n185 0.14
R8332 IREF.n202 IREF.n201 0.14
R8333 IREF.n211 IREF.n181 0.14
R8334 IREF.n212 IREF.n211 0.14
R8335 IREF.n213 IREF.n177 0.14
R8336 IREF.n221 IREF.n177 0.14
R8337 IREF.n228 IREF.n175 0.14
R8338 IREF.n229 IREF.n228 0.14
R8339 IREF.n230 IREF.n173 0.14
R8340 IREF.n234 IREF.n173 0.14
R8341 IREF.n395 IREF.n394 0.14
R8342 IREF.n394 IREF.n235 0.14
R8343 IREF.n387 IREF.n386 0.14
R8344 IREF.n386 IREF.n240 0.14
R8345 IREF.n379 IREF.n378 0.14
R8346 IREF.n378 IREF.n245 0.14
R8347 IREF.n371 IREF.n251 0.14
R8348 IREF.n371 IREF.n370 0.14
R8349 IREF.n362 IREF.n252 0.14
R8350 IREF.n362 IREF.n361 0.14
R8351 IREF.n353 IREF.n256 0.14
R8352 IREF.n353 IREF.n352 0.14
R8353 IREF.n344 IREF.n261 0.14
R8354 IREF.n344 IREF.n343 0.14
R8355 IREF.n268 IREF.n265 0.14
R8356 IREF.n334 IREF.n268 0.14
R8357 IREF.n329 IREF.n328 0.14
R8358 IREF.n328 IREF.n327 0.14
R8359 IREF.n323 IREF.n271 0.14
R8360 IREF.n323 IREF.n322 0.14
R8361 IREF.n321 IREF.n274 0.14
R8362 IREF.n314 IREF.n274 0.14
R8363 IREF.n313 IREF.n280 0.14
R8364 IREF.n306 IREF.n280 0.14
R8365 IREF.n305 IREF.n285 0.14
R8366 IREF.n298 IREF.n285 0.14
R8367 IREF.n297 IREF.n296 0.14
R8368 IREF.n197 IREF.n196 0.14
R8369 IREF.n197 IREF.n183 0.14
R8370 IREF.n206 IREF.n205 0.14
R8371 IREF.n206 IREF.n179 0.14
R8372 IREF.n217 IREF.n216 0.14
R8373 IREF.n217 IREF.n170 0.14
R8374 IREF.n397 IREF.n171 0.14
R8375 IREF.n391 IREF.n171 0.14
R8376 IREF.n390 IREF.n238 0.14
R8377 IREF.n383 IREF.n238 0.14
R8378 IREF.n382 IREF.n243 0.14
R8379 IREF.n375 IREF.n243 0.14
R8380 IREF.n374 IREF.n248 0.14
R8381 IREF.n368 IREF.n248 0.14
R8382 IREF.n367 IREF.n254 0.14
R8383 IREF.n258 IREF.n254 0.14
R8384 IREF.n358 IREF.n357 0.14
R8385 IREF.n357 IREF.n259 0.14
R8386 IREF.n349 IREF.n348 0.14
R8387 IREF.n348 IREF.n263 0.14
R8388 IREF.n339 IREF.n338 0.14
R8389 IREF.n338 IREF.n267 0.14
R8390 IREF.n318 IREF.n275 0.14
R8391 IREF.n318 IREF.n317 0.14
R8392 IREF.n310 IREF.n277 0.14
R8393 IREF.n310 IREF.n309 0.14
R8394 IREF.n302 IREF.n282 0.14
R8395 IREF.n302 IREF.n301 0.14
R8396 IREF.n293 IREF.n287 0.14
R8397 IREF.n418 IREF.n413 0.14
R8398 IREF.n426 IREF.n425 0.14
R8399 IREF.n427 IREF.n426 0.14
R8400 IREF.n434 IREF.n409 0.14
R8401 IREF.n435 IREF.n434 0.14
R8402 IREF.n436 IREF.n405 0.14
R8403 IREF.n442 IREF.n405 0.14
R8404 IREF.n449 IREF.n403 0.14
R8405 IREF.n450 IREF.n449 0.14
R8406 IREF.n451 IREF.n401 0.14
R8407 IREF.n455 IREF.n401 0.14
R8408 IREF.n457 IREF.n456 0.14
R8409 IREF.n456 IREF.n168 0.14
R8410 IREF.n466 IREF.n465 0.14
R8411 IREF.n466 IREF.n163 0.14
R8412 IREF.n473 IREF.n472 0.14
R8413 IREF.n475 IREF.n473 0.14
R8414 IREF.n474 IREF.n159 0.14
R8415 IREF.n483 IREF.n159 0.14
R8416 IREF.n485 IREF.n484 0.14
R8417 IREF.n484 IREF.n156 0.14
R8418 IREF.n494 IREF.n493 0.14
R8419 IREF.n494 IREF.n151 0.14
R8420 IREF.n501 IREF.n500 0.14
R8421 IREF.n503 IREF.n501 0.14
R8422 IREF.n502 IREF.n147 0.14
R8423 IREF.n511 IREF.n147 0.14
R8424 IREF.n518 IREF.n145 0.14
R8425 IREF.n519 IREF.n518 0.14
R8426 IREF.n520 IREF.n143 0.14
R8427 IREF.n524 IREF.n143 0.14
R8428 IREF.n526 IREF.n525 0.14
R8429 IREF.n527 IREF.n526 0.14
R8430 IREF.n532 IREF.n531 0.14
R8431 IREF.n533 IREF.n532 0.14
R8432 IREF.n537 IREF.n534 0.14
R8433 IREF.n538 IREF.n537 0.14
R8434 IREF.n542 IREF.n539 0.14
R8435 IREF.n421 IREF.n420 0.14
R8436 IREF.n423 IREF.n422 0.14
R8437 IREF.n422 IREF.n411 0.14
R8438 IREF.n432 IREF.n430 0.14
R8439 IREF.n432 IREF.n431 0.14
R8440 IREF.n439 IREF.n407 0.14
R8441 IREF.n440 IREF.n439 0.14
R8442 IREF.n461 IREF.n460 0.14
R8443 IREF.n462 IREF.n461 0.14
R8444 IREF.n468 IREF.n166 0.14
R8445 IREF.n469 IREF.n468 0.14
R8446 IREF.n470 IREF.n161 0.14
R8447 IREF.n477 IREF.n161 0.14
R8448 IREF.n479 IREF.n478 0.14
R8449 IREF.n479 IREF.n158 0.14
R8450 IREF.n489 IREF.n488 0.14
R8451 IREF.n490 IREF.n489 0.14
R8452 IREF.n496 IREF.n154 0.14
R8453 IREF.n497 IREF.n496 0.14
R8454 IREF.n498 IREF.n149 0.14
R8455 IREF.n505 IREF.n149 0.14
R8456 IREF.n507 IREF.n506 0.14
R8457 IREF.n507 IREF.n141 0.14
R8458 IREF.n561 IREF.n142 0.14
R8459 IREF.n556 IREF.n142 0.14
R8460 IREF.n555 IREF.n554 0.14
R8461 IREF.n554 IREF.n529 0.14
R8462 IREF.n550 IREF.n549 0.14
R8463 IREF.n549 IREF.n536 0.14
R8464 IREF.n545 IREF.n544 0.14
R8465 IREF.n614 IREF.n610 0.14
R8466 IREF.n623 IREF.n622 0.14
R8467 IREF.n623 IREF.n606 0.14
R8468 IREF.n633 IREF.n632 0.14
R8469 IREF.n634 IREF.n633 0.14
R8470 IREF.n642 IREF.n602 0.14
R8471 IREF.n659 IREF.n642 0.14
R8472 IREF.n654 IREF.n653 0.14
R8473 IREF.n653 IREF.n652 0.14
R8474 IREF.n648 IREF.n645 0.14
R8475 IREF.n648 IREF.n599 0.14
R8476 IREF.n667 IREF.n666 0.14
R8477 IREF.n667 IREF.n595 0.14
R8478 IREF.n676 IREF.n675 0.14
R8479 IREF.n676 IREF.n591 0.14
R8480 IREF.n686 IREF.n685 0.14
R8481 IREF.n687 IREF.n686 0.14
R8482 IREF.n695 IREF.n587 0.14
R8483 IREF.n696 IREF.n695 0.14
R8484 IREF.n704 IREF.n583 0.14
R8485 IREF.n705 IREF.n704 0.14
R8486 IREF.n713 IREF.n579 0.14
R8487 IREF.n714 IREF.n713 0.14
R8488 IREF.n723 IREF.n575 0.14
R8489 IREF.n724 IREF.n723 0.14
R8490 IREF.n725 IREF.n571 0.14
R8491 IREF.n733 IREF.n571 0.14
R8492 IREF.n740 IREF.n569 0.14
R8493 IREF.n741 IREF.n740 0.14
R8494 IREF.n742 IREF.n567 0.14
R8495 IREF.n746 IREF.n567 0.14
R8496 IREF.n790 IREF.n789 0.14
R8497 IREF.n789 IREF.n747 0.14
R8498 IREF.n782 IREF.n781 0.14
R8499 IREF.n781 IREF.n752 0.14
R8500 IREF.n774 IREF.n773 0.14
R8501 IREF.n773 IREF.n757 0.14
R8502 IREF.n766 IREF.n763 0.14
R8503 IREF.n618 IREF.n608 0.14
R8504 IREF.n626 IREF.n608 0.14
R8505 IREF.n627 IREF.n604 0.14
R8506 IREF.n637 IREF.n604 0.14
R8507 IREF.n638 IREF.n600 0.14
R8508 IREF.n661 IREF.n600 0.14
R8509 IREF.n663 IREF.n597 0.14
R8510 IREF.n670 IREF.n597 0.14
R8511 IREF.n671 IREF.n593 0.14
R8512 IREF.n679 IREF.n593 0.14
R8513 IREF.n680 IREF.n589 0.14
R8514 IREF.n690 IREF.n589 0.14
R8515 IREF.n691 IREF.n585 0.14
R8516 IREF.n698 IREF.n585 0.14
R8517 IREF.n700 IREF.n699 0.14
R8518 IREF.n700 IREF.n581 0.14
R8519 IREF.n709 IREF.n708 0.14
R8520 IREF.n709 IREF.n577 0.14
R8521 IREF.n718 IREF.n717 0.14
R8522 IREF.n718 IREF.n573 0.14
R8523 IREF.n729 IREF.n728 0.14
R8524 IREF.n729 IREF.n564 0.14
R8525 IREF.n792 IREF.n565 0.14
R8526 IREF.n786 IREF.n565 0.14
R8527 IREF.n785 IREF.n750 0.14
R8528 IREF.n778 IREF.n750 0.14
R8529 IREF.n777 IREF.n755 0.14
R8530 IREF.n770 IREF.n755 0.14
R8531 IREF.n769 IREF.n760 0.14
R8532 IREF.n71 IREF.n70 0.14
R8533 IREF.n77 IREF.n63 0.14
R8534 IREF.n78 IREF.n77 0.14
R8535 IREF.n79 IREF.n58 0.14
R8536 IREF.n86 IREF.n58 0.14
R8537 IREF.n88 IREF.n87 0.14
R8538 IREF.n88 IREF.n50 0.14
R8539 IREF.n1299 IREF.n51 0.14
R8540 IREF.n1294 IREF.n51 0.14
R8541 IREF.n1293 IREF.n1292 0.14
R8542 IREF.n1292 IREF.n110 0.14
R8543 IREF.n1288 IREF.n1287 0.14
R8544 IREF.n1287 IREF.n117 0.14
R8545 IREF.n1283 IREF.n1282 0.14
R8546 IREF.n1282 IREF.n1281 0.14
R8547 IREF.n1274 IREF.n122 0.14
R8548 IREF.n1274 IREF.n1273 0.14
R8549 IREF.n1272 IREF.n127 0.14
R8550 IREF.n1267 IREF.n127 0.14
R8551 IREF.n1266 IREF.n1265 0.14
R8552 IREF.n1265 IREF.n133 0.14
R8553 IREF.n1261 IREF.n1260 0.14
R8554 IREF.n1260 IREF.n1259 0.14
R8555 IREF.n1242 IREF.n1241 0.14
R8556 IREF.n1241 IREF.n1209 0.14
R8557 IREF.n1237 IREF.n1236 0.14
R8558 IREF.n1236 IREF.n1213 0.14
R8559 IREF.n1232 IREF.n1231 0.14
R8560 IREF.n1231 IREF.n1218 0.14
R8561 IREF.n1227 IREF.n1226 0.14
R8562 IREF.n881 IREF.n878 0.14
R8563 IREF.n887 IREF.n886 0.14
R8564 IREF.n888 IREF.n887 0.14
R8565 IREF.n892 IREF.n876 0.14
R8566 IREF.n893 IREF.n892 0.14
R8567 IREF.n900 IREF.n899 0.14
R8568 IREF.n900 IREF.n873 0.14
R8569 IREF.n906 IREF.n905 0.14
R8570 IREF.n907 IREF.n906 0.14
R8571 IREF.n912 IREF.n871 0.14
R8572 IREF.n913 IREF.n912 0.14
R8573 IREF.n914 IREF.n869 0.14
R8574 IREF.n918 IREF.n869 0.14
R8575 IREF.n921 IREF.n920 0.14
R8576 IREF.n922 IREF.n921 0.14
R8577 IREF.n927 IREF.n867 0.14
R8578 IREF.n928 IREF.n927 0.14
R8579 IREF.n929 IREF.n865 0.14
R8580 IREF.n934 IREF.n865 0.14
R8581 IREF.n936 IREF.n935 0.14
R8582 IREF.n936 IREF.n862 0.14
R8583 IREF.n959 IREF.n863 0.14
R8584 IREF.n954 IREF.n863 0.14
R8585 IREF.n953 IREF.n952 0.14
R8586 IREF.n952 IREF.n944 0.14
R8587 IREF.n835 IREF.n830 0.14
R8588 IREF.n840 IREF.n830 0.14
R8589 IREF.n842 IREF.n841 0.14
R8590 IREF.n842 IREF.n827 0.14
R8591 IREF.n1023 IREF.n828 0.14
R8592 IREF.n1018 IREF.n828 0.14
R8593 IREF.n1017 IREF.n1016 0.14
R8594 IREF.n1016 IREF.n850 0.14
R8595 IREF.n1011 IREF.n1010 0.14
R8596 IREF.n1010 IREF.n1009 0.14
R8597 IREF.n1005 IREF.n852 0.14
R8598 IREF.n1005 IREF.n1004 0.14
R8599 IREF.n999 IREF.n998 0.14
R8600 IREF.n998 IREF.n997 0.14
R8601 IREF.n993 IREF.n857 0.14
R8602 IREF.n993 IREF.n992 0.14
R8603 IREF.n988 IREF.n860 0.14
R8604 IREF.n988 IREF.n987 0.14
R8605 IREF.n981 IREF.n980 0.14
R8606 IREF.n980 IREF.n979 0.14
R8607 IREF.n975 IREF.n964 0.14
R8608 IREF.n975 IREF.n974 0.14
R8609 IREF.n970 IREF.n967 0.14
R8610 IREF.n1035 IREF.n1034 0.14
R8611 IREF.n1036 IREF.n1029 0.14
R8612 IREF.n1041 IREF.n1029 0.14
R8613 IREF.n1043 IREF.n1042 0.14
R8614 IREF.n1043 IREF.n1026 0.14
R8615 IREF.n1124 IREF.n1027 0.14
R8616 IREF.n1119 IREF.n1027 0.14
R8617 IREF.n1118 IREF.n1117 0.14
R8618 IREF.n1117 IREF.n1051 0.14
R8619 IREF.n1113 IREF.n1112 0.14
R8620 IREF.n1112 IREF.n1054 0.14
R8621 IREF.n1108 IREF.n1107 0.14
R8622 IREF.n1107 IREF.n1106 0.14
R8623 IREF.n1104 IREF.n1056 0.14
R8624 IREF.n1100 IREF.n1056 0.14
R8625 IREF.n1099 IREF.n1098 0.14
R8626 IREF.n1098 IREF.n1058 0.14
R8627 IREF.n1094 IREF.n1093 0.14
R8628 IREF.n1093 IREF.n1061 0.14
R8629 IREF.n1089 IREF.n1088 0.14
R8630 IREF.n1088 IREF.n1087 0.14
R8631 IREF.n1081 IREF.n1080 0.14
R8632 IREF.n1080 IREF.n1066 0.14
R8633 IREF.n1076 IREF.n1075 0.14
R8634 IREF.n1075 IREF.n1068 0.14
R8635 IREF.n820 IREF.n813 0.14
R8636 IREF.n821 IREF.n820 0.14
R8637 IREF.n825 IREF.n811 0.14
R8638 IREF.n1129 IREF.n825 0.14
R8639 IREF.n1136 IREF.n809 0.14
R8640 IREF.n1137 IREF.n1136 0.14
R8641 IREF.n1141 IREF.n807 0.14
R8642 IREF.n1142 IREF.n1141 0.14
R8643 IREF.n1147 IREF.n805 0.14
R8644 IREF.n1148 IREF.n1147 0.14
R8645 IREF.n1149 IREF.n803 0.14
R8646 IREF.n1153 IREF.n803 0.14
R8647 IREF.n1160 IREF.n801 0.14
R8648 IREF.n1161 IREF.n1160 0.14
R8649 IREF.n1162 IREF.n799 0.14
R8650 IREF.n1167 IREF.n799 0.14
R8651 IREF.n1169 IREF.n1168 0.14
R8652 IREF.n1169 IREF.n796 0.14
R8653 IREF.n1194 IREF.n797 0.14
R8654 IREF.n1189 IREF.n797 0.14
R8655 IREF.n1188 IREF.n1187 0.14
R8656 IREF.n1187 IREF.n1177 0.14
R8657 IREF.n1182 IREF.n1181 0.14
R8658 IREF.n1367 IREF.n1359 0.14
R8659 IREF.n1368 IREF.n1367 0.14
R8660 IREF.n1369 IREF.n1357 0.14
R8661 IREF.n1373 IREF.n1357 0.14
R8662 IREF.n1385 IREF.n1378 0.14
R8663 IREF.n1385 IREF.n1384 0.14
R8664 IREF.n7 IREF.n5 0.14
R8665 IREF.n12 IREF.n5 0.14
R8666 IREF.n13 IREF.n4 0.14
R8667 IREF.n16 IREF.n4 0.14
R8668 IREF.n17 IREF.n3 0.14
R8669 IREF.n21 IREF.n3 0.14
R8670 IREF.n1396 IREF.n22 0.14
R8671 IREF.n36 IREF.n35 0.1355
R8672 IREF.n1395 IREF.n23 0.1355
R8673 IREF.n1392 IREF.n1356 0.120905
R8674 IREF.n939 IREF.n938 0.118921
R8675 IREF.n894 IREF.n875 0.118921
R8676 IREF.n1086 IREF.n1064 0.118921
R8677 IREF.n1046 IREF.n1045 0.118921
R8678 IREF.n958 IREF.n957 0.116553
R8679 IREF.n898 IREF.n874 0.116553
R8680 IREF.n1082 IREF.n1065 0.116553
R8681 IREF.n1123 IREF.n1122 0.116553
R8682 IREF.n945 IREF.n943 0.114184
R8683 IREF.n925 IREF.n924 0.114184
R8684 IREF.n904 IREF.n903 0.114184
R8685 IREF.n1077 IREF.n1067 0.114184
R8686 IREF.n1059 IREF.n1057 0.114184
R8687 IREF.n1052 IREF.n1050 0.114184
R8688 IREF.n1254 IREF.n1253 0.109179
R8689 IREF.n1249 IREF.n1248 0.109179
R8690 IREF.n96 IREF.n95 0.109179
R8691 IREF.n102 IREF.n53 0.109179
R8692 IREF.n515 IREF.n514 0.109179
R8693 IREF.n521 IREF.n144 0.109179
R8694 IREF.n446 IREF.n445 0.109179
R8695 IREF.n452 IREF.n402 0.109179
R8696 IREF.n1234 IREF.n1233 0.107155
R8697 IREF.n1268 IREF.n132 0.107155
R8698 IREF.n1290 IREF.n1289 0.107155
R8699 IREF.n80 IREF.n61 0.107155
R8700 IREF.n552 IREF.n551 0.107155
R8701 IREF.n499 IREF.n152 0.107155
R8702 IREF.n471 IREF.n164 0.107155
R8703 IREF.n429 IREF.n428 0.107155
R8704 IREF.n1239 IREF.n1238 0.103632
R8705 IREF.n1271 IREF.n126 0.103632
R8706 IREF.n1295 IREF.n109 0.103632
R8707 IREF.n73 IREF.n72 0.103632
R8708 IREF.n557 IREF.n528 0.103632
R8709 IREF.n492 IREF.n491 0.103632
R8710 IREF.n464 IREF.n463 0.103632
R8711 IREF.n424 IREF.n414 0.103632
R8712 IREF.n331 IREF.n330 0.102991
R8713 IREF.n326 IREF.n325 0.102991
R8714 IREF.n225 IREF.n224 0.102991
R8715 IREF.n231 IREF.n174 0.102991
R8716 IREF.n737 IREF.n736 0.102991
R8717 IREF.n743 IREF.n568 0.102991
R8718 IREF.n656 IREF.n655 0.102991
R8719 IREF.n651 IREF.n650 0.102991
R8720 IREF.n949 IREF.n946 0.0987895
R8721 IREF.n931 IREF.n930 0.0987895
R8722 IREF.n910 IREF.n909 0.0987895
R8723 IREF.n885 IREF.n884 0.0987895
R8724 IREF.n1072 IREF.n1069 0.0987895
R8725 IREF.n1095 IREF.n1060 0.0987895
R8726 IREF.n1114 IREF.n1053 0.0987895
R8727 IREF.n1038 IREF.n1037 0.0987895
R8728 IREF.n315 IREF.n279 0.0933826
R8729 IREF.n360 IREF.n359 0.0933826
R8730 IREF.n389 IREF.n237 0.0933826
R8731 IREF.n195 IREF.n194 0.0933826
R8732 IREF.n784 IREF.n749 0.0933826
R8733 IREF.n707 IREF.n706 0.0933826
R8734 IREF.n672 IREF.n596 0.0933826
R8735 IREF.n619 IREF.n611 0.0933826
R8736 IREF.n307 IREF.n284 0.092742
R8737 IREF.n351 IREF.n350 0.092742
R8738 IREF.n381 IREF.n242 0.092742
R8739 IREF.n204 IREF.n203 0.092742
R8740 IREF.n776 IREF.n754 0.092742
R8741 IREF.n716 IREF.n715 0.092742
R8742 IREF.n681 IREF.n592 0.092742
R8743 IREF.n628 IREF.n607 0.092742
R8744 IREF IREF.n1397 0.0822105
R8745 IREF.n1229 IREF.n1228 0.0821726
R8746 IREF.n1263 IREF.n1262 0.0821726
R8747 IREF.n1285 IREF.n1284 0.0821726
R8748 IREF.n85 IREF.n57 0.0821726
R8749 IREF.n299 IREF.n289 0.0821726
R8750 IREF.n342 IREF.n341 0.0821726
R8751 IREF.n249 IREF.n247 0.0821726
R8752 IREF.n214 IREF.n180 0.0821726
R8753 IREF.n547 IREF.n546 0.0821726
R8754 IREF.n504 IREF.n148 0.0821726
R8755 IREF.n476 IREF.n160 0.0821726
R8756 IREF.n437 IREF.n408 0.0821726
R8757 IREF.n761 IREF.n759 0.0821726
R8758 IREF.n726 IREF.n574 0.0821726
R8759 IREF.n688 IREF.n588 0.0821726
R8760 IREF.n635 IREF.n603 0.0821726
R8761 IREF.n36 IREF.n31 0.0733942
R8762 IREF.n932 IREF.n931 0.0490526
R8763 IREF.n911 IREF.n910 0.0490526
R8764 IREF.n884 IREF.n877 0.0490526
R8765 IREF.n1092 IREF.n1060 0.0490526
R8766 IREF.n1111 IREF.n1053 0.0490526
R8767 IREF.n1039 IREF.n1038 0.0490526
R8768 IREF.n1253 IREF.n1203 0.0426132
R8769 IREF.n1248 IREF.n1247 0.0426132
R8770 IREF.n98 IREF.n96 0.0426132
R8771 IREF.n103 IREF.n102 0.0426132
R8772 IREF.n517 IREF.n515 0.0426132
R8773 IREF.n522 IREF.n521 0.0426132
R8774 IREF.n448 IREF.n446 0.0426132
R8775 IREF.n453 IREF.n452 0.0426132
R8776 IREF.n1255 IREF.n1254 0.0412547
R8777 IREF.n1249 IREF.n1205 0.0412547
R8778 IREF.n95 IREF.n55 0.0412547
R8779 IREF.n97 IREF.n53 0.0412547
R8780 IREF.n514 IREF.n146 0.0412547
R8781 IREF.n516 IREF.n144 0.0412547
R8782 IREF.n445 IREF.n404 0.0412547
R8783 IREF.n447 IREF.n402 0.0412547
R8784 IREF.n1240 IREF.n1239 0.0402153
R8785 IREF.n1235 IREF.n1234 0.0402153
R8786 IREF.n1230 IREF.n1229 0.0402153
R8787 IREF.n1228 IREF.n1222 0.0402153
R8788 IREF.n1275 IREF.n126 0.0402153
R8789 IREF.n1269 IREF.n1268 0.0402153
R8790 IREF.n1264 IREF.n1263 0.0402153
R8791 IREF.n1262 IREF.n139 0.0402153
R8792 IREF.n1296 IREF.n1295 0.0402153
R8793 IREF.n1291 IREF.n1290 0.0402153
R8794 IREF.n1286 IREF.n1285 0.0402153
R8795 IREF.n1284 IREF.n121 0.0402153
R8796 IREF.n72 IREF.n66 0.0402153
R8797 IREF.n76 IREF.n61 0.0402153
R8798 IREF.n85 IREF.n59 0.0402153
R8799 IREF.n89 IREF.n57 0.0402153
R8800 IREF.n330 IREF.n270 0.0402153
R8801 IREF.n325 IREF.n324 0.0402153
R8802 IREF.n227 IREF.n225 0.0402153
R8803 IREF.n232 IREF.n231 0.0402153
R8804 IREF.n558 IREF.n557 0.0402153
R8805 IREF.n553 IREF.n552 0.0402153
R8806 IREF.n548 IREF.n547 0.0402153
R8807 IREF.n546 IREF.n540 0.0402153
R8808 IREF.n491 IREF.n157 0.0402153
R8809 IREF.n495 IREF.n152 0.0402153
R8810 IREF.n504 IREF.n150 0.0402153
R8811 IREF.n508 IREF.n148 0.0402153
R8812 IREF.n463 IREF.n169 0.0402153
R8813 IREF.n467 IREF.n164 0.0402153
R8814 IREF.n476 IREF.n162 0.0402153
R8815 IREF.n480 IREF.n160 0.0402153
R8816 IREF.n419 IREF.n414 0.0402153
R8817 IREF.n428 IREF.n412 0.0402153
R8818 IREF.n433 IREF.n408 0.0402153
R8819 IREF.n438 IREF.n437 0.0402153
R8820 IREF.n739 IREF.n737 0.0402153
R8821 IREF.n744 IREF.n743 0.0402153
R8822 IREF.n655 IREF.n644 0.0402153
R8823 IREF.n650 IREF.n649 0.0402153
R8824 IREF.n332 IREF.n331 0.0389342
R8825 IREF.n326 IREF.n272 0.0389342
R8826 IREF.n224 IREF.n176 0.0389342
R8827 IREF.n226 IREF.n174 0.0389342
R8828 IREF.n736 IREF.n570 0.0389342
R8829 IREF.n738 IREF.n568 0.0389342
R8830 IREF.n657 IREF.n656 0.0389342
R8831 IREF.n651 IREF.n646 0.0389342
R8832 IREF.n295 IREF.n291 0.0338096
R8833 IREF.n340 IREF.n266 0.0338096
R8834 IREF.n373 IREF.n372 0.0338096
R8835 IREF.n215 IREF.n178 0.0338096
R8836 IREF.n768 IREF.n767 0.0338096
R8837 IREF.n727 IREF.n572 0.0338096
R8838 IREF.n694 IREF.n692 0.0338096
R8839 IREF.n641 IREF.n639 0.0338096
R8840 IREF.n951 IREF.n945 0.0336579
R8841 IREF.n926 IREF.n925 0.0336579
R8842 IREF.n903 IREF.n872 0.0336579
R8843 IREF.n882 IREF.n879 0.0336579
R8844 IREF.n1074 IREF.n1067 0.0336579
R8845 IREF.n1097 IREF.n1059 0.0336579
R8846 IREF.n1116 IREF.n1052 0.0336579
R8847 IREF.n1033 IREF.n1032 0.0336579
R8848 IREF.n1225 IREF.n1223 0.0325285
R8849 IREF.n1258 IREF.n1200 0.0325285
R8850 IREF.n1280 IREF.n123 0.0325285
R8851 IREF.n91 IREF.n90 0.0325285
R8852 IREF.n292 IREF.n290 0.0325285
R8853 IREF.n336 IREF.n335 0.0325285
R8854 IREF.n369 IREF.n253 0.0325285
R8855 IREF.n220 IREF.n219 0.0325285
R8856 IREF.n543 IREF.n541 0.0325285
R8857 IREF.n510 IREF.n509 0.0325285
R8858 IREF.n482 IREF.n481 0.0325285
R8859 IREF.n441 IREF.n406 0.0325285
R8860 IREF.n765 IREF.n764 0.0325285
R8861 IREF.n732 IREF.n731 0.0325285
R8862 IREF.n697 IREF.n586 0.0325285
R8863 IREF.n660 IREF.n601 0.0325285
R8864 IREF.n1243 IREF.n1208 0.0318879
R8865 IREF.n1277 IREF.n1276 0.0318879
R8866 IREF.n1298 IREF.n1297 0.0318879
R8867 IREF.n69 IREF.n68 0.0318879
R8868 IREF.n560 IREF.n559 0.0318879
R8869 IREF.n487 IREF.n486 0.0318879
R8870 IREF.n459 IREF.n458 0.0318879
R8871 IREF.n417 IREF.n416 0.0318879
R8872 IREF.n957 IREF.n956 0.0312895
R8873 IREF.n919 IREF.n868 0.0312895
R8874 IREF.n901 IREF.n874 0.0312895
R8875 IREF.n1079 IREF.n1065 0.0312895
R8876 IREF.n1103 IREF.n1102 0.0312895
R8877 IREF.n1122 IREF.n1121 0.0312895
R8878 IREF.n1238 IREF.n1212 0.0312473
R8879 IREF.n1271 IREF.n1270 0.0312473
R8880 IREF.n111 IREF.n109 0.0312473
R8881 IREF.n73 IREF.n64 0.0312473
R8882 IREF.n530 IREF.n528 0.0312473
R8883 IREF.n492 IREF.n155 0.0312473
R8884 IREF.n464 IREF.n167 0.0312473
R8885 IREF.n424 IREF.n415 0.0312473
R8886 IREF.n320 IREF.n319 0.0306068
R8887 IREF.n316 IREF.n278 0.0306068
R8888 IREF.n366 IREF.n365 0.0306068
R8889 IREF.n363 IREF.n255 0.0306068
R8890 IREF.n396 IREF.n172 0.0306068
R8891 IREF.n393 IREF.n392 0.0306068
R8892 IREF.n191 IREF.n188 0.0306068
R8893 IREF.n791 IREF.n566 0.0306068
R8894 IREF.n788 IREF.n787 0.0306068
R8895 IREF.n701 IREF.n584 0.0306068
R8896 IREF.n703 IREF.n582 0.0306068
R8897 IREF.n665 IREF.n664 0.0306068
R8898 IREF.n669 IREF.n668 0.0306068
R8899 IREF.n616 IREF.n615 0.0306068
R8900 IREF.n312 IREF.n311 0.0299662
R8901 IREF.n308 IREF.n283 0.0299662
R8902 IREF.n356 IREF.n257 0.0299662
R8903 IREF.n354 IREF.n260 0.0299662
R8904 IREF.n388 IREF.n239 0.0299662
R8905 IREF.n385 IREF.n384 0.0299662
R8906 IREF.n198 IREF.n186 0.0299662
R8907 IREF.n200 IREF.n184 0.0299662
R8908 IREF.n783 IREF.n751 0.0299662
R8909 IREF.n780 IREF.n779 0.0299662
R8910 IREF.n710 IREF.n580 0.0299662
R8911 IREF.n712 IREF.n578 0.0299662
R8912 IREF.n674 IREF.n673 0.0299662
R8913 IREF.n678 IREF.n677 0.0299662
R8914 IREF.n621 IREF.n620 0.0299662
R8915 IREF.n625 IREF.n624 0.0299662
R8916 IREF.n938 IREF.n937 0.0289211
R8917 IREF.n917 IREF.n916 0.0289211
R8918 IREF.n891 IREF.n875 0.0289211
R8919 IREF.n1064 IREF.n1062 0.0289211
R8920 IREF.n1105 IREF.n1055 0.0289211
R8921 IREF.n1045 IREF.n1044 0.0289211
R8922 IREF.n1233 IREF.n1217 0.0270836
R8923 IREF.n134 IREF.n132 0.0270836
R8924 IREF.n1289 IREF.n116 0.0270836
R8925 IREF.n80 IREF.n62 0.0270836
R8926 IREF.n551 IREF.n535 0.0270836
R8927 IREF.n499 IREF.n153 0.0270836
R8928 IREF.n471 IREF.n165 0.0270836
R8929 IREF.n429 IREF.n410 0.0270836
R8930 IREF.n304 IREF.n303 0.0258025
R8931 IREF.n300 IREF.n288 0.0258025
R8932 IREF.n347 IREF.n262 0.0258025
R8933 IREF.n345 IREF.n264 0.0258025
R8934 IREF.n380 IREF.n244 0.0258025
R8935 IREF.n377 IREF.n376 0.0258025
R8936 IREF.n207 IREF.n182 0.0258025
R8937 IREF.n210 IREF.n209 0.0258025
R8938 IREF.n775 IREF.n756 0.0258025
R8939 IREF.n772 IREF.n771 0.0258025
R8940 IREF.n719 IREF.n576 0.0258025
R8941 IREF.n722 IREF.n721 0.0258025
R8942 IREF.n684 IREF.n683 0.0258025
R8943 IREF.n689 IREF.n590 0.0258025
R8944 IREF.n631 IREF.n630 0.0258025
R8945 IREF.n636 IREF.n605 0.0258025
R8946 IREF.n190 IREF.n189 0.0170406
R8947 IREF.n613 IREF.n612 0.0170406
R8948 IREF.n304 IREF.n284 0.0149128
R8949 IREF.n300 IREF.n299 0.0149128
R8950 IREF.n350 IREF.n262 0.0149128
R8951 IREF.n342 IREF.n264 0.0149128
R8952 IREF.n381 IREF.n380 0.0149128
R8953 IREF.n376 IREF.n247 0.0149128
R8954 IREF.n204 IREF.n182 0.0149128
R8955 IREF.n209 IREF.n180 0.0149128
R8956 IREF.n776 IREF.n775 0.0149128
R8957 IREF.n771 IREF.n759 0.0149128
R8958 IREF.n716 IREF.n576 0.0149128
R8959 IREF.n721 IREF.n574 0.0149128
R8960 IREF.n684 IREF.n681 0.0149128
R8961 IREF.n689 IREF.n688 0.0149128
R8962 IREF.n631 IREF.n628 0.0149128
R8963 IREF.n636 IREF.n635 0.0149128
R8964 IREF.n1230 IREF.n1217 0.0136317
R8965 IREF.n1264 IREF.n134 0.0136317
R8966 IREF.n1286 IREF.n116 0.0136317
R8967 IREF.n62 IREF.n59 0.0136317
R8968 IREF.n288 IREF.n286 0.0136317
R8969 IREF.n346 IREF.n345 0.0136317
R8970 IREF.n377 IREF.n246 0.0136317
R8971 IREF.n210 IREF.n208 0.0136317
R8972 IREF.n548 IREF.n535 0.0136317
R8973 IREF.n153 IREF.n150 0.0136317
R8974 IREF.n165 IREF.n162 0.0136317
R8975 IREF.n433 IREF.n410 0.0136317
R8976 IREF.n772 IREF.n758 0.0136317
R8977 IREF.n722 IREF.n720 0.0136317
R8978 IREF.n682 IREF.n590 0.0136317
R8979 IREF.n629 IREF.n605 0.0136317
R8980 IREF.n312 IREF.n279 0.0107491
R8981 IREF.n308 IREF.n307 0.0107491
R8982 IREF.n359 IREF.n257 0.0107491
R8983 IREF.n351 IREF.n260 0.0107491
R8984 IREF.n389 IREF.n388 0.0107491
R8985 IREF.n384 IREF.n242 0.0107491
R8986 IREF.n195 IREF.n186 0.0107491
R8987 IREF.n203 IREF.n184 0.0107491
R8988 IREF.n784 IREF.n783 0.0107491
R8989 IREF.n779 IREF.n754 0.0107491
R8990 IREF.n707 IREF.n580 0.0107491
R8991 IREF.n715 IREF.n578 0.0107491
R8992 IREF.n674 IREF.n672 0.0107491
R8993 IREF.n678 IREF.n592 0.0107491
R8994 IREF.n621 IREF.n619 0.0107491
R8995 IREF.n625 IREF.n607 0.0107491
R8996 IREF.n316 IREF.n315 0.0101085
R8997 IREF.n360 IREF.n255 0.0101085
R8998 IREF.n392 IREF.n237 0.0101085
R8999 IREF.n194 IREF.n188 0.0101085
R9000 IREF.n787 IREF.n749 0.0101085
R9001 IREF.n706 IREF.n582 0.0101085
R9002 IREF.n669 IREF.n596 0.0101085
R9003 IREF.n616 IREF.n611 0.0101085
R9004 IREF.n1235 IREF.n1212 0.00946797
R9005 IREF.n1270 IREF.n1269 0.00946797
R9006 IREF.n1291 IREF.n111 0.00946797
R9007 IREF.n76 IREF.n64 0.00946797
R9008 IREF.n283 IREF.n281 0.00946797
R9009 IREF.n355 IREF.n354 0.00946797
R9010 IREF.n385 IREF.n241 0.00946797
R9011 IREF.n200 IREF.n199 0.00946797
R9012 IREF.n553 IREF.n530 0.00946797
R9013 IREF.n495 IREF.n155 0.00946797
R9014 IREF.n467 IREF.n167 0.00946797
R9015 IREF.n415 IREF.n412 0.00946797
R9016 IREF.n780 IREF.n753 0.00946797
R9017 IREF.n712 IREF.n711 0.00946797
R9018 IREF.n677 IREF.n594 0.00946797
R9019 IREF.n624 IREF.n609 0.00946797
R9020 IREF.n1240 IREF.n1208 0.0088274
R9021 IREF.n1276 IREF.n1275 0.0088274
R9022 IREF.n1297 IREF.n1296 0.0088274
R9023 IREF.n68 IREF.n66 0.0088274
R9024 IREF.n278 IREF.n276 0.0088274
R9025 IREF.n364 IREF.n363 0.0088274
R9026 IREF.n393 IREF.n236 0.0088274
R9027 IREF.n191 IREF.n190 0.0088274
R9028 IREF.n559 IREF.n558 0.0088274
R9029 IREF.n486 IREF.n157 0.0088274
R9030 IREF.n458 IREF.n169 0.0088274
R9031 IREF.n419 IREF.n417 0.0088274
R9032 IREF.n788 IREF.n748 0.0088274
R9033 IREF.n703 IREF.n702 0.0088274
R9034 IREF.n668 IREF.n598 0.0088274
R9035 IREF.n615 IREF.n613 0.0088274
R9036 IREF.n1223 IREF.n1222 0.00818683
R9037 IREF.n1200 IREF.n139 0.00818683
R9038 IREF.n123 IREF.n121 0.00818683
R9039 IREF.n90 IREF.n89 0.00818683
R9040 IREF.n541 IREF.n540 0.00818683
R9041 IREF.n509 IREF.n508 0.00818683
R9042 IREF.n481 IREF.n480 0.00818683
R9043 IREF.n438 IREF.n406 0.00818683
R9044 IREF.n291 IREF.n289 0.00690569
R9045 IREF.n295 IREF.n294 0.00690569
R9046 IREF.n341 IREF.n340 0.00690569
R9047 IREF.n337 IREF.n266 0.00690569
R9048 IREF.n373 IREF.n249 0.00690569
R9049 IREF.n372 IREF.n250 0.00690569
R9050 IREF.n215 IREF.n214 0.00690569
R9051 IREF.n218 IREF.n178 0.00690569
R9052 IREF.n768 IREF.n761 0.00690569
R9053 IREF.n767 IREF.n762 0.00690569
R9054 IREF.n727 IREF.n726 0.00690569
R9055 IREF.n730 IREF.n572 0.00690569
R9056 IREF.n692 IREF.n588 0.00690569
R9057 IREF.n694 IREF.n693 0.00690569
R9058 IREF.n639 IREF.n603 0.00690569
R9059 IREF.n641 IREF.n640 0.00690569
R9060 IREF.n1192 IREF.n1191 0.00523684
R9061 IREF.n1186 IREF.n1185 0.00523684
R9062 IREF.n1179 IREF.n1178 0.00523684
R9063 IREF.n1159 IREF.n1158 0.00523684
R9064 IREF.n1165 IREF.n1164 0.00523684
R9065 IREF.n1171 IREF.n1170 0.00523684
R9066 IREF.n1135 IREF.n808 0.00523684
R9067 IREF.n1140 IREF.n806 0.00523684
R9068 IREF.n1146 IREF.n1145 0.00523684
R9069 IREF.n1152 IREF.n1151 0.00523684
R9070 IREF.n819 IREF.n812 0.00523684
R9071 IREF.n824 IREF.n810 0.00523684
R9072 IREF.n965 IREF.n963 0.00523684
R9073 IREF.n976 IREF.n966 0.00523684
R9074 IREF.n971 IREF.n968 0.00523684
R9075 IREF.n858 IREF.n856 0.00523684
R9076 IREF.n994 IREF.n859 0.00523684
R9077 IREF.n989 IREF.n861 0.00523684
R9078 IREF.n1021 IREF.n1020 0.00523684
R9079 IREF.n1015 IREF.n1014 0.00523684
R9080 IREF.n853 IREF.n851 0.00523684
R9081 IREF.n1006 IREF.n854 0.00523684
R9082 IREF.n838 IREF.n837 0.00523684
R9083 IREF.n844 IREF.n843 0.00523684
R9084 IREF.n1366 IREF.n1365 0.00523684
R9085 IREF.n1372 IREF.n1371 0.00523684
R9086 IREF.n1396 IREF.n1395 0.005
R9087 IREF.n1205 IREF.n1203 0.00185849
R9088 IREF.n1247 IREF.n1206 0.00185849
R9089 IREF.n98 IREF.n97 0.00185849
R9090 IREF.n104 IREF.n103 0.00185849
R9091 IREF.n517 IREF.n516 0.00185849
R9092 IREF.n523 IREF.n522 0.00185849
R9093 IREF.n448 IREF.n447 0.00185849
R9094 IREF.n454 IREF.n453 0.00185849
R9095 IREF.n319 IREF.n276 0.00178114
R9096 IREF.n311 IREF.n281 0.00178114
R9097 IREF.n303 IREF.n286 0.00178114
R9098 IREF.n294 IREF.n292 0.00178114
R9099 IREF.n365 IREF.n364 0.00178114
R9100 IREF.n356 IREF.n355 0.00178114
R9101 IREF.n347 IREF.n346 0.00178114
R9102 IREF.n337 IREF.n336 0.00178114
R9103 IREF.n236 IREF.n172 0.00178114
R9104 IREF.n241 IREF.n239 0.00178114
R9105 IREF.n246 IREF.n244 0.00178114
R9106 IREF.n253 IREF.n250 0.00178114
R9107 IREF.n272 IREF.n270 0.00178114
R9108 IREF.n324 IREF.n273 0.00178114
R9109 IREF.n227 IREF.n226 0.00178114
R9110 IREF.n233 IREF.n232 0.00178114
R9111 IREF.n199 IREF.n198 0.00178114
R9112 IREF.n208 IREF.n207 0.00178114
R9113 IREF.n219 IREF.n218 0.00178114
R9114 IREF.n748 IREF.n566 0.00178114
R9115 IREF.n753 IREF.n751 0.00178114
R9116 IREF.n758 IREF.n756 0.00178114
R9117 IREF.n764 IREF.n762 0.00178114
R9118 IREF.n702 IREF.n701 0.00178114
R9119 IREF.n711 IREF.n710 0.00178114
R9120 IREF.n720 IREF.n719 0.00178114
R9121 IREF.n731 IREF.n730 0.00178114
R9122 IREF.n664 IREF.n598 0.00178114
R9123 IREF.n673 IREF.n594 0.00178114
R9124 IREF.n683 IREF.n682 0.00178114
R9125 IREF.n693 IREF.n586 0.00178114
R9126 IREF.n739 IREF.n738 0.00178114
R9127 IREF.n745 IREF.n744 0.00178114
R9128 IREF.n646 IREF.n644 0.00178114
R9129 IREF.n649 IREF.n647 0.00178114
R9130 IREF.n620 IREF.n609 0.00178114
R9131 IREF.n630 IREF.n629 0.00178114
R9132 IREF.n640 IREF.n601 0.00178114
R9133 IREF.n45 IREF.n44 0.00168421
R9134 IREF.n20 IREF.n19 0.00168421
R9135 IREF.n15 IREF.n14 0.00168421
R9136 IREF.n11 IREF.n10 0.00168421
R9137 IREF.n1397 IREF.n2 0.00168421
R9138 a_n11737_n15980.n137 a_n11737_n15980.n136 12.734
R9139 a_n11737_n15980.n63 a_n11737_n15980.t27 8.41809
R9140 a_n11737_n15980.n64 a_n11737_n15980.t36 8.41809
R9141 a_n11737_n15980.n63 a_n11737_n15980.t44 8.37125
R9142 a_n11737_n15980.n67 a_n11737_n15980.t63 8.37125
R9143 a_n11737_n15980.n64 a_n11737_n15980.t48 8.37125
R9144 a_n11737_n15980.n110 a_n11737_n15980.t29 8.33806
R9145 a_n11737_n15980.n104 a_n11737_n15980.t62 8.3366
R9146 a_n11737_n15980.n89 a_n11737_n15980.t56 8.26493
R9147 a_n11737_n15980.n123 a_n11737_n15980.t39 8.2602
R9148 a_n11737_n15980.n17 a_n11737_n15980.t35 8.06917
R9149 a_n11737_n15980.n28 a_n11737_n15980.t42 8.06917
R9150 a_n11737_n15980.n13 a_n11737_n15980.t28 8.06917
R9151 a_n11737_n15980.n13 a_n11737_n15980.t41 8.06917
R9152 a_n11737_n15980.n11 a_n11737_n15980.t53 8.06917
R9153 a_n11737_n15980.n11 a_n11737_n15980.t40 8.06917
R9154 a_n11737_n15980.n69 a_n11737_n15980.t52 8.06917
R9155 a_n11737_n15980.n17 a_n11737_n15980.t64 8.06917
R9156 a_n11737_n15980.n30 a_n11737_n15980.t34 8.06917
R9157 a_n11737_n15980.n7 a_n11737_n15980.t50 8.06917
R9158 a_n11737_n15980.n7 a_n11737_n15980.t37 8.06917
R9159 a_n11737_n15980.n32 a_n11737_n15980.t49 8.06917
R9160 a_n11737_n15980.n83 a_n11737_n15980.t55 8.06917
R9161 a_n11737_n15980.n3 a_n11737_n15980.t45 8.06917
R9162 a_n11737_n15980.n3 a_n11737_n15980.t54 8.06917
R9163 a_n11737_n15980.n21 a_n11737_n15980.t26 8.06917
R9164 a_n11737_n15980.n21 a_n11737_n15980.t58 8.06917
R9165 a_n11737_n15980.n77 a_n11737_n15980.t25 8.06917
R9166 a_n11737_n15980.n103 a_n11737_n15980.t51 8.06917
R9167 a_n11737_n15980.n0 a_n11737_n15980.t61 8.06917
R9168 a_n11737_n15980.n101 a_n11737_n15980.t32 8.06917
R9169 a_n11737_n15980.n100 a_n11737_n15980.t60 8.06917
R9170 a_n11737_n15980.n99 a_n11737_n15980.t31 8.06917
R9171 a_n11737_n15980.n97 a_n11737_n15980.t57 8.06917
R9172 a_n11737_n15980.n90 a_n11737_n15980.t43 8.06917
R9173 a_n11737_n15980.n117 a_n11737_n15980.t30 8.06917
R9174 a_n11737_n15980.n111 a_n11737_n15980.t59 8.06917
R9175 a_n11737_n15980.n119 a_n11737_n15980.t46 8.06917
R9176 a_n11737_n15980.n120 a_n11737_n15980.t33 8.06917
R9177 a_n11737_n15980.n121 a_n11737_n15980.t47 8.06917
R9178 a_n11737_n15980.n124 a_n11737_n15980.t24 8.06917
R9179 a_n11737_n15980.n130 a_n11737_n15980.t38 8.06917
R9180 a_n11737_n15980.n66 a_n11737_n15980.t0 6.65728
R9181 a_n11737_n15980.n49 a_n11737_n15980.t13 6.51495
R9182 a_n11737_n15980.n140 a_n11737_n15980.n42 6.40828
R9183 a_n11737_n15980.n44 a_n11737_n15980.n43 6.37877
R9184 a_n11737_n15980.n66 a_n11737_n15980.t1 5.74368
R9185 a_n11737_n15980.n51 a_n11737_n15980.n50 5.24318
R9186 a_n11737_n15980.n71 a_n11737_n15980.n31 2.4223
R9187 a_n11737_n15980.n78 a_n11737_n15980.n33 2.42484
R9188 a_n11737_n15980.n79 a_n11737_n15980.n33 2.4256
R9189 a_n11737_n15980.n39 a_n11737_n15980.n38 2.24636
R9190 a_n11737_n15980.t12 a_n11737_n15980.n35 5.26436
R9191 a_n11737_n15980.n60 a_n11737_n15980.n44 4.60825
R9192 a_n11737_n15980.n34 a_n11737_n15980.n151 3.79435
R9193 a_n11737_n15980.n38 a_n11737_n15980.n140 4.59811
R9194 a_n11737_n15980.n22 a_n11737_n15980.n21 0.592766
R9195 a_n11737_n15980.n12 a_n11737_n15980.n11 0.592803
R9196 a_n11737_n15980.n15 a_n11737_n15980.n13 0.591918
R9197 a_n11737_n15980.n17 a_n11737_n15980.n18 0.591826
R9198 a_n11737_n15980.n37 a_n11737_n15980.n36 2.24389
R9199 a_n11737_n15980.n55 a_n11737_n15980.n45 4.5005
R9200 a_n11737_n15980.n10 a_n11737_n15980.n73 4.5005
R9201 a_n11737_n15980.n13 a_n11737_n15980.n14 0.591264
R9202 a_n11737_n15980.n74 a_n11737_n15980.n24 4.5005
R9203 a_n11737_n15980.n31 a_n11737_n15980.n30 0.0133501
R9204 a_n11737_n15980.n16 a_n11737_n15980.n71 4.5005
R9205 a_n11737_n15980.n19 a_n11737_n15980.n17 0.604195
R9206 a_n11737_n15980.n29 a_n11737_n15980.n70 4.5005
R9207 a_n11737_n15980.n76 a_n11737_n15980.n75 4.5005
R9208 a_n11737_n15980.n28 a_n11737_n15980.n27 0.0143905
R9209 a_n11737_n15980.n20 a_n11737_n15980.n81 4.5005
R9210 a_n11737_n15980.n2 a_n11737_n15980.n82 4.5005
R9211 a_n11737_n15980.n3 a_n11737_n15980.n4 0.591675
R9212 a_n11737_n15980.n9 a_n11737_n15980.n7 0.604671
R9213 a_n11737_n15980.n6 a_n11737_n15980.n78 4.5005
R9214 a_n11737_n15980.n32 a_n11737_n15980.n33 0.0107891
R9215 a_n11737_n15980.n7 a_n11737_n15980.n8 0.604671
R9216 a_n11737_n15980.n79 a_n11737_n15980.n6 4.5005
R9217 a_n11737_n15980.n2 a_n11737_n15980.n23 4.5005
R9218 a_n11737_n15980.n5 a_n11737_n15980.n3 0.591675
R9219 a_n11737_n15980.n91 a_n11737_n15980.n88 4.5005
R9220 a_n11737_n15980.n93 a_n11737_n15980.n92 4.5005
R9221 a_n11737_n15980.n94 a_n11737_n15980.n87 4.5005
R9222 a_n11737_n15980.n96 a_n11737_n15980.n95 4.5005
R9223 a_n11737_n15980.n98 a_n11737_n15980.n86 4.5005
R9224 a_n11737_n15980.n1 a_n11737_n15980.n0 1.44113
R9225 a_n11737_n15980.n105 a_n11737_n15980.n102 4.5005
R9226 a_n11737_n15980.n118 a_n11737_n15980.n107 4.5005
R9227 a_n11737_n15980.n116 a_n11737_n15980.n115 4.5005
R9228 a_n11737_n15980.n114 a_n11737_n15980.n109 4.5005
R9229 a_n11737_n15980.n113 a_n11737_n15980.n112 4.5005
R9230 a_n11737_n15980.n133 a_n11737_n15980.n132 4.5005
R9231 a_n11737_n15980.n131 a_n11737_n15980.n108 4.5005
R9232 a_n11737_n15980.n129 a_n11737_n15980.n128 4.5005
R9233 a_n11737_n15980.n127 a_n11737_n15980.n122 4.5005
R9234 a_n11737_n15980.n126 a_n11737_n15980.n125 4.5005
R9235 a_n11737_n15980.n149 a_n11737_n15980.n148 4.5005
R9236 a_n11737_n15980.n40 a_n11737_n15980.n41 2.23676
R9237 a_n11737_n15980.n36 a_n11737_n15980.n46 3.79594
R9238 a_n11737_n15980.n152 a_n11737_n15980.n40 3.79475
R9239 a_n11737_n15980.n147 a_n11737_n15980.t19 3.77936
R9240 a_n11737_n15980.n56 a_n11737_n15980.t5 3.77818
R9241 a_n11737_n15980.n49 a_n11737_n15980.n48 3.77318
R9242 a_n11737_n15980.n145 a_n11737_n15980.n144 3.77081
R9243 a_n11737_n15980.n54 a_n11737_n15980.n53 3.75571
R9244 a_n11737_n15980.n138 a_n11737_n15980.n62 2.69513
R9245 a_n11737_n15980.n84 a_n11737_n15980.n82 2.4256
R9246 a_n11737_n15980.n23 a_n11737_n15980.n84 2.42484
R9247 a_n11737_n15980.n31 a_n11737_n15980.n70 2.43326
R9248 a_n11737_n15980.n38 a_n11737_n15980.n142 2.32949
R9249 a_n11737_n15980.n135 a_n11737_n15980.n106 2.30989
R9250 a_n11737_n15980.n60 a_n11737_n15980.n59 2.30818
R9251 a_n11737_n15980.n147 a_n11737_n15980.n146 2.24481
R9252 a_n11737_n15980.n61 a_n11737_n15980.n60 2.2442
R9253 a_n11737_n15980.n57 a_n11737_n15980.n56 2.24358
R9254 a_n11737_n15980.n80 a_n11737_n15980.n77 2.23529
R9255 a_n11737_n15980.n72 a_n11737_n15980.n69 2.23423
R9256 a_n11737_n15980.n106 a_n11737_n15980.n86 2.18975
R9257 a_n11737_n15980.n134 a_n11737_n15980.n107 2.16725
R9258 a_n11737_n15980.n26 a_n11737_n15980.n5 2.4981
R9259 a_n11737_n15980.n136 a_n11737_n15980.n85 2.07557
R9260 a_n11737_n15980.n85 a_n11737_n15980.n25 2.07182
R9261 a_n11737_n15980.n25 a_n11737_n15980.n15 2.4644
R9262 a_n11737_n15980.n67 a_n11737_n15980.n66 1.7613
R9263 a_n11737_n15980.n65 a_n11737_n15980.n63 1.55888
R9264 a_n11737_n15980.n85 a_n11737_n15980.n26 1.5005
R9265 a_n11737_n15980.n135 a_n11737_n15980.n134 1.5005
R9266 a_n11737_n15980.n65 a_n11737_n15980.n64 1.5005
R9267 a_n11737_n15980.n68 a_n11737_n15980.n67 1.5005
R9268 a_n11737_n15980.n139 a_n11737_n15980.n138 1.5005
R9269 a_n11737_n15980.n151 a_n11737_n15980.t8 1.4705
R9270 a_n11737_n15980.n151 a_n11737_n15980.n150 1.4705
R9271 a_n11737_n15980.n53 a_n11737_n15980.t3 1.4705
R9272 a_n11737_n15980.n53 a_n11737_n15980.n52 1.4705
R9273 a_n11737_n15980.n48 a_n11737_n15980.t18 1.4705
R9274 a_n11737_n15980.n48 a_n11737_n15980.n47 1.4705
R9275 a_n11737_n15980.n59 a_n11737_n15980.t10 1.4705
R9276 a_n11737_n15980.n59 a_n11737_n15980.n58 1.4705
R9277 a_n11737_n15980.n142 a_n11737_n15980.t17 1.4705
R9278 a_n11737_n15980.n142 a_n11737_n15980.n141 1.4705
R9279 a_n11737_n15980.n144 a_n11737_n15980.t4 1.4705
R9280 a_n11737_n15980.n144 a_n11737_n15980.n143 1.4705
R9281 a_n11737_n15980.n89 a_n11737_n15980.n88 1.39514
R9282 a_n11737_n15980.n126 a_n11737_n15980.n123 1.39105
R9283 a_n11737_n15980.n136 a_n11737_n15980.n135 1.35453
R9284 a_n11737_n15980.n51 a_n11737_n15980.n49 1.27228
R9285 a_n11737_n15980.n99 a_n11737_n15980.n98 1.26997
R9286 a_n11737_n15980.n0 a_n11737_n15980.n101 1.24392
R9287 a_n11737_n15980.n119 a_n11737_n15980.n118 1.24204
R9288 a_n11737_n15980.n146 a_n11737_n15980.n145 1.20603
R9289 a_n11737_n15980.n132 a_n11737_n15980.n121 1.20414
R9290 a_n11737_n15980.n105 a_n11737_n15980.n104 1.14132
R9291 a_n11737_n15980.n61 a_n11737_n15980.n57 1.13952
R9292 a_n11737_n15980.n113 a_n11737_n15980.n110 1.13598
R9293 a_n11737_n15980.n37 a_n11737_n15980.n54 1.20574
R9294 a_n11737_n15980.n41 a_n11737_n15980.n34 1.24017
R9295 a_n11737_n15980.n138 a_n11737_n15980.n137 0.963743
R9296 a_n11737_n15980.n54 a_n11737_n15980.n51 0.937067
R9297 a_n11737_n15980.n106 a_n11737_n15980.n1 0.888471
R9298 a_n11737_n15980.n134 a_n11737_n15980.n133 0.71825
R9299 a_n11737_n15980.n100 a_n11737_n15980.n99 0.663658
R9300 a_n11737_n15980.n101 a_n11737_n15980.n100 0.663658
R9301 a_n11737_n15980.n121 a_n11737_n15980.n120 0.655156
R9302 a_n11737_n15980.n120 a_n11737_n15980.n119 0.655156
R9303 a_n11737_n15980.n124 a_n11737_n15980.n123 0.439529
R9304 a_n11737_n15980.n90 a_n11737_n15980.n89 0.432797
R9305 a_n11737_n15980.n129 a_n11737_n15980.n122 0.379447
R9306 a_n11737_n15980.n112 a_n11737_n15980.n109 0.379447
R9307 a_n11737_n15980.n71 a_n11737_n15980.n19 0.745981
R9308 a_n11737_n15980.n9 a_n11737_n15980.n78 0.745252
R9309 a_n11737_n15980.n8 a_n11737_n15980.n79 0.745252
R9310 a_n11737_n15980.n1 a_n11737_n15980.n105 0.498861
R9311 a_n11737_n15980.n73 a_n11737_n15980.n12 0.756573
R9312 a_n11737_n15980.n18 a_n11737_n15980.n70 0.756388
R9313 a_n11737_n15980.n15 a_n11737_n15980.n76 0.756711
R9314 a_n11737_n15980.n81 a_n11737_n15980.n22 0.756011
R9315 a_n11737_n15980.n114 a_n11737_n15980.n113 0.3605
R9316 a_n11737_n15980.n128 a_n11737_n15980.n127 0.3605
R9317 a_n11737_n15980.n104 a_n11737_n15980.n103 0.335806
R9318 a_n11737_n15980.n111 a_n11737_n15980.n110 0.33475
R9319 a_n11737_n15980.n92 a_n11737_n15980.n87 0.302474
R9320 a_n11737_n15980.n94 a_n11737_n15980.n93 0.287375
R9321 a_n11737_n15980.n137 a_n11737_n15980.n68 0.277797
R9322 a_n11737_n15980.n73 a_n11737_n15980.n72 0.208888
R9323 a_n11737_n15980.n81 a_n11737_n15980.n80 0.20887
R9324 a_n11737_n15980.n57 a_n11737_n15980.n45 0.208394
R9325 a_n11737_n15980.n149 a_n11737_n15980.n146 0.208357
R9326 a_n11737_n15980.n68 a_n11737_n15980.n65 0.168946
R9327 a_n11737_n15980.n37 a_n11737_n15980.n45 0.233116
R9328 a_n11737_n15980.n92 a_n11737_n15980.n91 0.147342
R9329 a_n11737_n15980.n96 a_n11737_n15980.n87 0.147342
R9330 a_n11737_n15980.n132 a_n11737_n15980.n131 0.147342
R9331 a_n11737_n15980.n125 a_n11737_n15980.n122 0.147342
R9332 a_n11737_n15980.n116 a_n11737_n15980.n109 0.147342
R9333 a_n11737_n15980.n41 a_n11737_n15980.n149 0.211956
R9334 a_n11737_n15980.n148 a_n11737_n15980.n40 0.142388
R9335 a_n11737_n15980.n62 a_n11737_n15980.n44 0.14
R9336 a_n11737_n15980.n72 a_n11737_n15980.n19 1.12746
R9337 a_n11737_n15980.n14 a_n11737_n15980.n12 1.49123
R9338 a_n11737_n15980.n14 a_n11737_n15980.n24 0.772202
R9339 a_n11737_n15980.n18 a_n11737_n15980.n25 1.21369
R9340 a_n11737_n15980.n76 a_n11737_n15980.n27 2.42126
R9341 a_n11737_n15980.n80 a_n11737_n15980.n9 1.12837
R9342 a_n11737_n15980.n4 a_n11737_n15980.n22 1.49118
R9343 a_n11737_n15980.n82 a_n11737_n15980.n4 0.772883
R9344 a_n11737_n15980.n8 a_n11737_n15980.n26 1.21186
R9345 a_n11737_n15980.n5 a_n11737_n15980.n23 0.772883
R9346 a_n11737_n15980.n93 a_n11737_n15980.n88 0.14
R9347 a_n11737_n15980.n95 a_n11737_n15980.n94 0.14
R9348 a_n11737_n15980.n95 a_n11737_n15980.n86 0.14
R9349 a_n11737_n15980.n115 a_n11737_n15980.n114 0.14
R9350 a_n11737_n15980.n115 a_n11737_n15980.n107 0.14
R9351 a_n11737_n15980.n133 a_n11737_n15980.n108 0.14
R9352 a_n11737_n15980.n128 a_n11737_n15980.n108 0.14
R9353 a_n11737_n15980.n127 a_n11737_n15980.n126 0.14
R9354 a_n11737_n15980.n35 a_n11737_n15980.n39 1.19679
R9355 a_n11737_n15980.n145 a_n11737_n15980.n35 0.932624
R9356 a_n11737_n15980.t20 a_n11737_n15980.n34 6.53226
R9357 a_n11737_n15980.n118 a_n11737_n15980.n117 0.137868
R9358 a_n11737_n15980.n55 a_n11737_n15980.n36 0.137318
R9359 a_n11737_n15980.n140 a_n11737_n15980.n139 0.131
R9360 a_n11737_n15980.n103 a_n11737_n15980.n102 0.128395
R9361 a_n11737_n15980.n112 a_n11737_n15980.n111 0.128395
R9362 a_n11737_n15980.n130 a_n11737_n15980.n129 0.118921
R9363 a_n11737_n15980.n98 a_n11737_n15980.n97 0.114184
R9364 a_n11737_n15980.n56 a_n11737_n15980.n55 0.110782
R9365 a_n11737_n15980.n148 a_n11737_n15980.n147 0.105711
R9366 a_n11737_n15980.n62 a_n11737_n15980.n61 0.0688756
R9367 a_n11737_n15980.n32 a_n11737_n15980.n6 0.0402153
R9368 a_n11737_n15980.n91 a_n11737_n15980.n90 0.0348421
R9369 a_n11737_n15980.n20 a_n11737_n15980.n77 0.0344623
R9370 a_n11737_n15980.n97 a_n11737_n15980.n96 0.0336579
R9371 a_n11737_n15980.n10 a_n11737_n15980.n69 0.0325285
R9372 a_n11737_n15980.n30 a_n11737_n15980.n29 0.0299662
R9373 a_n11737_n15980.n131 a_n11737_n15980.n130 0.0289211
R9374 a_n11737_n15980.n2 a_n11737_n15980.n83 0.0283648
R9375 a_n11737_n15980.n74 a_n11737_n15980.n28 0.0258025
R9376 a_n11737_n15980.n84 a_n11737_n15980.n83 0.0226397
R9377 a_n11737_n15980.n125 a_n11737_n15980.n124 0.0194474
R9378 a_n11737_n15980.n75 a_n11737_n15980.n74 0.0149128
R9379 a_n11737_n15980.n16 a_n11737_n15980.n29 0.0107491
R9380 a_n11737_n15980.n117 a_n11737_n15980.n116 0.00997368
R9381 a_n11737_n15980.n139 a_n11737_n15980.n39 0.0777922
R9382 a_n11737_n15980.n24 a_n11737_n15980.n27 2.43637
R9383 a_n11737_n15980.n0 a_n11737_n15980.n102 0.6755
R9384 a_n11737_n15980.n3 a_n11737_n15980.n2 0.369148
R9385 a_n11737_n15980.n75 a_n11737_n15980.n13 0.354735
R9386 a_n11737_n15980.n7 a_n11737_n15980.n6 0.347689
R9387 a_n11737_n15980.n17 a_n11737_n15980.n16 0.347689
R9388 a_n11737_n15980.n21 a_n11737_n15980.n20 0.346915
R9389 a_n11737_n15980.n11 a_n11737_n15980.n10 0.32719
R9390 a_n13990_8177.n72 a_n13990_8177.n69 7.94229
R9391 a_n13990_8177.n140 a_n13990_8177.n135 7.94229
R9392 a_n13990_8177.n359 a_n13990_8177.n355 7.22198
R9393 a_n13990_8177.n417 a_n13990_8177.n416 7.22198
R9394 a_n13990_8177.n337 a_n13990_8177.n334 6.77653
R9395 a_n13990_8177.n314 a_n13990_8177.n311 6.77653
R9396 a_n13990_8177.n323 a_n13990_8177.t266 6.7761
R9397 a_n13990_8177.n320 a_n13990_8177.t164 6.7761
R9398 a_n13990_8177.n21 a_n13990_8177.n306 6.77231
R9399 a_n13990_8177.n31 a_n13990_8177.n367 6.77231
R9400 a_n13990_8177.n300 a_n13990_8177.t44 6.58663
R9401 a_n13990_8177.n238 a_n13990_8177.t64 6.58663
R9402 a_n13990_8177.n515 a_n13990_8177.n514 6.50088
R9403 a_n13990_8177.n471 a_n13990_8177.n470 6.50088
R9404 a_n13990_8177.n301 a_n13990_8177.n297 5.95439
R9405 a_n13990_8177.n239 a_n13990_8177.n235 5.95439
R9406 a_n13990_8177.n68 a_n13990_8177.n67 5.69423
R9407 a_n13990_8177.n74 a_n13990_8177.n73 5.69423
R9408 a_n13990_8177.n139 a_n13990_8177.n138 5.69423
R9409 a_n13990_8177.n132 a_n13990_8177.n131 5.69423
R9410 a_n13990_8177.n343 a_n13990_8177.t231 5.50607
R9411 a_n13990_8177.n338 a_n13990_8177.t195 5.50607
R9412 a_n13990_8177.n386 a_n13990_8177.t129 5.50607
R9413 a_n13990_8177.n315 a_n13990_8177.t264 5.50607
R9414 a_n13990_8177.n342 a_n13990_8177.n341 5.50475
R9415 a_n13990_8177.n348 a_n13990_8177.n347 5.50475
R9416 a_n13990_8177.n349 a_n13990_8177.t144 5.50475
R9417 a_n13990_8177.n340 a_n13990_8177.n339 5.50475
R9418 a_n13990_8177.n385 a_n13990_8177.n384 5.50475
R9419 a_n13990_8177.n391 a_n13990_8177.n390 5.50475
R9420 a_n13990_8177.n392 a_n13990_8177.t222 5.50475
R9421 a_n13990_8177.n317 a_n13990_8177.n316 5.50475
R9422 a_n13990_8177.n68 a_n13990_8177.n66 5.49558
R9423 a_n13990_8177.n139 a_n13990_8177.n137 5.49558
R9424 a_n13990_8177.n297 a_n13990_8177.t19 5.31528
R9425 a_n13990_8177.n235 a_n13990_8177.t6 5.31528
R9426 a_n13990_8177.n521 a_n13990_8177.n518 4.92758
R9427 a_n13990_8177.n432 a_n13990_8177.n429 4.92758
R9428 a_n13990_8177.n38 a_n13990_8177.n489 4.92217
R9429 a_n13990_8177.n45 a_n13990_8177.n440 4.92217
R9430 a_n13990_8177.n0 a_n13990_8177.n128 4.22068
R9431 a_n13990_8177.t157 a_n13990_8177.n1 5.69068
R9432 a_n13990_8177.n126 a_n13990_8177.n2 4.22068
R9433 a_n13990_8177.n3 a_n13990_8177.n63 4.22068
R9434 a_n13990_8177.n4 a_n13990_8177.t143 5.69068
R9435 a_n13990_8177.n5 a_n13990_8177.n61 4.22068
R9436 a_n13990_8177.n7 a_n13990_8177.n181 3.84173
R9437 a_n13990_8177.n10 a_n13990_8177.n171 3.84173
R9438 a_n13990_8177.n504 a_n13990_8177.n32 3.65107
R9439 a_n13990_8177.n502 a_n13990_8177.n33 3.65107
R9440 a_n13990_8177.n500 a_n13990_8177.n34 3.65107
R9441 a_n13990_8177.n498 a_n13990_8177.n35 3.65107
R9442 a_n13990_8177.n495 a_n13990_8177.n36 3.65107
R9443 a_n13990_8177.n493 a_n13990_8177.n37 3.65107
R9444 a_n13990_8177.n491 a_n13990_8177.n38 3.65107
R9445 a_n13990_8177.n39 a_n13990_8177.n454 3.65107
R9446 a_n13990_8177.n40 a_n13990_8177.n452 3.65107
R9447 a_n13990_8177.n41 a_n13990_8177.n450 3.65107
R9448 a_n13990_8177.n42 a_n13990_8177.n448 3.65107
R9449 a_n13990_8177.n446 a_n13990_8177.n43 3.65107
R9450 a_n13990_8177.n444 a_n13990_8177.n44 3.65107
R9451 a_n13990_8177.n442 a_n13990_8177.n45 3.65107
R9452 a_n13990_8177.n12 a_n13990_8177.n553 4.0312
R9453 a_n13990_8177.n551 a_n13990_8177.n13 5.5012
R9454 a_n13990_8177.t200 a_n13990_8177.n14 5.5012
R9455 a_n13990_8177.n550 a_n13990_8177.n15 4.0312
R9456 a_n13990_8177.n548 a_n13990_8177.n16 5.5012
R9457 a_n13990_8177.t165 a_n13990_8177.n17 5.5012
R9458 a_n13990_8177.n547 a_n13990_8177.n18 4.0312
R9459 a_n13990_8177.n309 a_n13990_8177.n19 5.5012
R9460 a_n13990_8177.t263 a_n13990_8177.n20 5.5012
R9461 a_n13990_8177.n308 a_n13990_8177.n21 4.0312
R9462 a_n13990_8177.n22 a_n13990_8177.n379 4.0312
R9463 a_n13990_8177.n377 a_n13990_8177.n23 5.5012
R9464 a_n13990_8177.t257 a_n13990_8177.n24 5.5012
R9465 a_n13990_8177.n376 a_n13990_8177.n25 4.0312
R9466 a_n13990_8177.n374 a_n13990_8177.n26 5.5012
R9467 a_n13990_8177.t169 a_n13990_8177.n27 5.5012
R9468 a_n13990_8177.n373 a_n13990_8177.n28 4.0312
R9469 a_n13990_8177.n370 a_n13990_8177.n29 5.5012
R9470 a_n13990_8177.t218 a_n13990_8177.n30 5.5012
R9471 a_n13990_8177.n369 a_n13990_8177.n31 4.0312
R9472 a_n13990_8177.n6 a_n13990_8177.n175 5.31173
R9473 a_n13990_8177.n8 a_n13990_8177.n179 5.31173
R9474 a_n13990_8177.n9 a_n13990_8177.n172 5.31173
R9475 a_n13990_8177.n11 a_n13990_8177.n169 5.31173
R9476 a_n13990_8177.n296 a_n13990_8177.n293 4.50663
R9477 a_n13990_8177.n234 a_n13990_8177.n168 4.50663
R9478 a_n13990_8177.n182 a_n13990_8177.n8 4.46113
R9479 a_n13990_8177.n358 a_n13990_8177.n357 4.24002
R9480 a_n13990_8177.n327 a_n13990_8177.n326 4.24002
R9481 a_n13990_8177.n415 a_n13990_8177.n414 4.24002
R9482 a_n13990_8177.n400 a_n13990_8177.n399 4.24002
R9483 a_n13990_8177.n72 a_n13990_8177.n71 4.22423
R9484 a_n13990_8177.n135 a_n13990_8177.n134 4.22423
R9485 a_n13990_8177.n463 a_n13990_8177.t286 4.06712
R9486 a_n13990_8177.n461 a_n13990_8177.t74 4.06712
R9487 a_n13990_8177.n507 a_n13990_8177.t337 4.06712
R9488 a_n13990_8177.n425 a_n13990_8177.t344 4.06712
R9489 a_n13990_8177.n152 a_n13990_8177.t114 4.05054
R9490 a_n13990_8177.n161 a_n13990_8177.n160 4.05054
R9491 a_n13990_8177.n163 a_n13990_8177.t214 4.05054
R9492 a_n13990_8177.n144 a_n13990_8177.n143 4.05054
R9493 a_n13990_8177.n47 a_n13990_8177.t181 4.05054
R9494 a_n13990_8177.n567 a_n13990_8177.n566 4.05054
R9495 a_n13990_8177.n563 a_n13990_8177.t106 4.05054
R9496 a_n13990_8177.n51 a_n13990_8177.n50 4.05054
R9497 a_n13990_8177.n84 a_n13990_8177.t260 4.05054
R9498 a_n13990_8177.n93 a_n13990_8177.n92 4.05054
R9499 a_n13990_8177.n95 a_n13990_8177.t228 4.05054
R9500 a_n13990_8177.n106 a_n13990_8177.n105 4.05054
R9501 a_n13990_8177.n108 a_n13990_8177.t140 4.05054
R9502 a_n13990_8177.n118 a_n13990_8177.n117 4.05054
R9503 a_n13990_8177.n120 a_n13990_8177.t188 4.05054
R9504 a_n13990_8177.n77 a_n13990_8177.n76 4.05054
R9505 a_n13990_8177.n323 a_n13990_8177.n322 4.03475
R9506 a_n13990_8177.n346 a_n13990_8177.n345 4.03475
R9507 a_n13990_8177.n352 a_n13990_8177.n351 4.03475
R9508 a_n13990_8177.n337 a_n13990_8177.n336 4.03475
R9509 a_n13990_8177.n320 a_n13990_8177.n319 4.03475
R9510 a_n13990_8177.n389 a_n13990_8177.n388 4.03475
R9511 a_n13990_8177.n395 a_n13990_8177.n394 4.03475
R9512 a_n13990_8177.n314 a_n13990_8177.n313 4.03475
R9513 a_n13990_8177.n508 a_n13990_8177.n506 3.96014
R9514 a_n13990_8177.n464 a_n13990_8177.n427 3.96014
R9515 a_n13990_8177.n152 a_n13990_8177.t145 3.87765
R9516 a_n13990_8177.n161 a_n13990_8177.n159 3.87765
R9517 a_n13990_8177.n163 a_n13990_8177.t116 3.87765
R9518 a_n13990_8177.n144 a_n13990_8177.n142 3.87765
R9519 a_n13990_8177.n47 a_n13990_8177.t209 3.87765
R9520 a_n13990_8177.n567 a_n13990_8177.n565 3.87765
R9521 a_n13990_8177.n563 a_n13990_8177.t244 3.87765
R9522 a_n13990_8177.n51 a_n13990_8177.n49 3.87765
R9523 a_n13990_8177.n84 a_n13990_8177.t247 3.87765
R9524 a_n13990_8177.n93 a_n13990_8177.n91 3.87765
R9525 a_n13990_8177.n95 a_n13990_8177.t223 3.87765
R9526 a_n13990_8177.n106 a_n13990_8177.n104 3.87765
R9527 a_n13990_8177.n108 a_n13990_8177.t128 3.87765
R9528 a_n13990_8177.n118 a_n13990_8177.n116 3.87765
R9529 a_n13990_8177.n120 a_n13990_8177.t179 3.87765
R9530 a_n13990_8177.n77 a_n13990_8177.n75 3.87765
R9531 a_n13990_8177.n463 a_n13990_8177.t288 3.86107
R9532 a_n13990_8177.n461 a_n13990_8177.t75 3.86107
R9533 a_n13990_8177.n507 a_n13990_8177.t284 3.86107
R9534 a_n13990_8177.n425 a_n13990_8177.t342 3.86107
R9535 a_n13990_8177.n300 a_n13990_8177.n299 3.84528
R9536 a_n13990_8177.n296 a_n13990_8177.n295 3.84528
R9537 a_n13990_8177.n238 a_n13990_8177.n237 3.84528
R9538 a_n13990_8177.n234 a_n13990_8177.n233 3.84528
R9539 a_n13990_8177.n285 a_n13990_8177.n279 3.79678
R9540 a_n13990_8177.n260 a_n13990_8177.n254 3.79678
R9541 a_n13990_8177.n200 a_n13990_8177.n194 3.79678
R9542 a_n13990_8177.n223 a_n13990_8177.n217 3.79678
R9543 a_n13990_8177.n524 a_n13990_8177.n521 3.79678
R9544 a_n13990_8177.n536 a_n13990_8177.n533 3.79678
R9545 a_n13990_8177.n435 a_n13990_8177.n432 3.79678
R9546 a_n13990_8177.n483 a_n13990_8177.n480 3.79678
R9547 a_n13990_8177.n243 a_n13990_8177.n11 3.87644
R9548 a_n13990_8177.n273 a_n13990_8177.n267 3.73034
R9549 a_n13990_8177.n230 a_n13990_8177.n206 3.73034
R9550 a_n13990_8177.n358 a_n13990_8177.n356 3.68818
R9551 a_n13990_8177.n327 a_n13990_8177.n325 3.68818
R9552 a_n13990_8177.n415 a_n13990_8177.n413 3.68818
R9553 a_n13990_8177.n400 a_n13990_8177.n398 3.68818
R9554 a_n13990_8177.n530 a_n13990_8177.n529 3.65581
R9555 a_n13990_8177.n533 a_n13990_8177.n532 3.65581
R9556 a_n13990_8177.n536 a_n13990_8177.n535 3.65581
R9557 a_n13990_8177.n539 a_n13990_8177.n538 3.65581
R9558 a_n13990_8177.n527 a_n13990_8177.n526 3.65581
R9559 a_n13990_8177.n524 a_n13990_8177.n523 3.65581
R9560 a_n13990_8177.n521 a_n13990_8177.n520 3.65581
R9561 a_n13990_8177.n486 a_n13990_8177.n485 3.65581
R9562 a_n13990_8177.n483 a_n13990_8177.n482 3.65581
R9563 a_n13990_8177.n480 a_n13990_8177.n479 3.65581
R9564 a_n13990_8177.n477 a_n13990_8177.n476 3.65581
R9565 a_n13990_8177.n438 a_n13990_8177.n437 3.65581
R9566 a_n13990_8177.n435 a_n13990_8177.n434 3.65581
R9567 a_n13990_8177.n432 a_n13990_8177.n431 3.65581
R9568 a_n13990_8177.n540 a_n13990_8177.n539 3.64443
R9569 a_n13990_8177.n477 a_n13990_8177.n474 3.64443
R9570 a_n13990_8177.n35 a_n13990_8177.n496 3.64223
R9571 a_n13990_8177.n455 a_n13990_8177.n42 3.64223
R9572 a_n13990_8177.n123 a_n13990_8177.n74 3.25667
R9573 a_n13990_8177.n366 a_n13990_8177.n365 3.23904
R9574 a_n13990_8177.n412 a_n13990_8177.n305 3.23904
R9575 a_n13990_8177.n2 a_n13990_8177.n124 3.15553
R9576 a_n13990_8177.n560 a_n13990_8177.n5 3.15553
R9577 a_n13990_8177.n301 a_n13990_8177.n300 3.00663
R9578 a_n13990_8177.n239 a_n13990_8177.n238 3.00663
R9579 a_n13990_8177.n248 a_n13990_8177.n245 2.7866
R9580 a_n13990_8177.n253 a_n13990_8177.n250 2.7866
R9581 a_n13990_8177.n259 a_n13990_8177.n256 2.7866
R9582 a_n13990_8177.n265 a_n13990_8177.n262 2.7866
R9583 a_n13990_8177.n272 a_n13990_8177.n269 2.7866
R9584 a_n13990_8177.n278 a_n13990_8177.n275 2.7866
R9585 a_n13990_8177.n284 a_n13990_8177.n281 2.7866
R9586 a_n13990_8177.n290 a_n13990_8177.n287 2.7866
R9587 a_n13990_8177.n211 a_n13990_8177.n208 2.7866
R9588 a_n13990_8177.n216 a_n13990_8177.n213 2.7866
R9589 a_n13990_8177.n222 a_n13990_8177.n219 2.7866
R9590 a_n13990_8177.n228 a_n13990_8177.n225 2.7866
R9591 a_n13990_8177.n205 a_n13990_8177.n202 2.7866
R9592 a_n13990_8177.n199 a_n13990_8177.n196 2.7866
R9593 a_n13990_8177.n193 a_n13990_8177.n190 2.7866
R9594 a_n13990_8177.n187 a_n13990_8177.n184 2.7866
R9595 a_n13990_8177.n364 a_n13990_8177.n363 2.77002
R9596 a_n13990_8177.n332 a_n13990_8177.n331 2.77002
R9597 a_n13990_8177.n411 a_n13990_8177.n410 2.77002
R9598 a_n13990_8177.n405 a_n13990_8177.n404 2.77002
R9599 a_n13990_8177.n83 a_n13990_8177.n77 2.73714
R9600 a_n13990_8177.n333 a_n13990_8177.n327 2.73714
R9601 a_n13990_8177.n406 a_n13990_8177.n400 2.73714
R9602 a_n13990_8177.n426 a_n13990_8177.n424 2.73714
R9603 a_n13990_8177.n462 a_n13990_8177.n460 2.73714
R9604 a_n13990_8177.n57 a_n13990_8177.n51 2.73714
R9605 a_n13990_8177.n158 a_n13990_8177.n152 2.73672
R9606 a_n13990_8177.n90 a_n13990_8177.n84 2.73672
R9607 a_n13990_8177.n254 a_n13990_8177.n248 2.73672
R9608 a_n13990_8177.n217 a_n13990_8177.n211 2.73672
R9609 a_n13990_8177.n109 a_n13990_8177.n107 2.60203
R9610 a_n13990_8177.n349 a_n13990_8177.n348 2.60203
R9611 a_n13990_8177.n392 a_n13990_8177.n391 2.60203
R9612 a_n13990_8177.n145 a_n13990_8177.n48 2.60203
R9613 a_n13990_8177.n469 a_n13990_8177.n466 2.59712
R9614 a_n13990_8177.n460 a_n13990_8177.n457 2.59712
R9615 a_n13990_8177.n513 a_n13990_8177.n510 2.59712
R9616 a_n13990_8177.n424 a_n13990_8177.n421 2.59712
R9617 a_n13990_8177.n157 a_n13990_8177.n156 2.58054
R9618 a_n13990_8177.n150 a_n13990_8177.n149 2.58054
R9619 a_n13990_8177.n56 a_n13990_8177.n55 2.58054
R9620 a_n13990_8177.n89 a_n13990_8177.n88 2.58054
R9621 a_n13990_8177.n102 a_n13990_8177.n101 2.58054
R9622 a_n13990_8177.n114 a_n13990_8177.n113 2.58054
R9623 a_n13990_8177.n82 a_n13990_8177.n81 2.58054
R9624 a_n13990_8177.n573 a_n13990_8177.n572 2.58054
R9625 a_n13990_8177.n121 a_n13990_8177.n119 2.53418
R9626 a_n13990_8177.n96 a_n13990_8177.n94 2.53418
R9627 a_n13990_8177.n568 a_n13990_8177.n564 2.53418
R9628 a_n13990_8177.n164 a_n13990_8177.n162 2.53418
R9629 a_n13990_8177.n340 a_n13990_8177.n338 2.52436
R9630 a_n13990_8177.n343 a_n13990_8177.n342 2.52436
R9631 a_n13990_8177.n317 a_n13990_8177.n315 2.52436
R9632 a_n13990_8177.n386 a_n13990_8177.n385 2.52436
R9633 a_n13990_8177.n132 a_n13990_8177.n58 2.51873
R9634 a_n13990_8177.n515 a_n13990_8177.n426 2.46014
R9635 a_n13990_8177.n471 a_n13990_8177.n462 2.46014
R9636 a_n13990_8177.n157 a_n13990_8177.n154 2.40765
R9637 a_n13990_8177.n150 a_n13990_8177.n147 2.40765
R9638 a_n13990_8177.n56 a_n13990_8177.n53 2.40765
R9639 a_n13990_8177.n89 a_n13990_8177.n86 2.40765
R9640 a_n13990_8177.n102 a_n13990_8177.n99 2.40765
R9641 a_n13990_8177.n114 a_n13990_8177.n111 2.40765
R9642 a_n13990_8177.n82 a_n13990_8177.n79 2.40765
R9643 a_n13990_8177.n572 a_n13990_8177.n571 2.40765
R9644 a_n13990_8177.n469 a_n13990_8177.n468 2.39107
R9645 a_n13990_8177.n460 a_n13990_8177.n459 2.39107
R9646 a_n13990_8177.n513 a_n13990_8177.n512 2.39107
R9647 a_n13990_8177.n424 a_n13990_8177.n423 2.39107
R9648 a_n13990_8177.n242 a_n13990_8177.n9 2.37644
R9649 a_n13990_8177.n178 a_n13990_8177.n6 2.37644
R9650 a_n13990_8177.n69 a_n13990_8177.n64 2.23844
R9651 a_n13990_8177.n364 a_n13990_8177.n361 2.21818
R9652 a_n13990_8177.n332 a_n13990_8177.n329 2.21818
R9653 a_n13990_8177.n411 a_n13990_8177.n408 2.21818
R9654 a_n13990_8177.n405 a_n13990_8177.n402 2.21818
R9655 a_n13990_8177.n248 a_n13990_8177.n247 2.2016
R9656 a_n13990_8177.n253 a_n13990_8177.n252 2.2016
R9657 a_n13990_8177.n259 a_n13990_8177.n258 2.2016
R9658 a_n13990_8177.n265 a_n13990_8177.n264 2.2016
R9659 a_n13990_8177.n272 a_n13990_8177.n271 2.2016
R9660 a_n13990_8177.n278 a_n13990_8177.n277 2.2016
R9661 a_n13990_8177.n284 a_n13990_8177.n283 2.2016
R9662 a_n13990_8177.n290 a_n13990_8177.n289 2.2016
R9663 a_n13990_8177.n211 a_n13990_8177.n210 2.2016
R9664 a_n13990_8177.n216 a_n13990_8177.n215 2.2016
R9665 a_n13990_8177.n222 a_n13990_8177.n221 2.2016
R9666 a_n13990_8177.n228 a_n13990_8177.n227 2.2016
R9667 a_n13990_8177.n205 a_n13990_8177.n204 2.2016
R9668 a_n13990_8177.n199 a_n13990_8177.n198 2.2016
R9669 a_n13990_8177.n193 a_n13990_8177.n192 2.2016
R9670 a_n13990_8177.n187 a_n13990_8177.n186 2.2016
R9671 a_n13990_8177.n354 a_n13990_8177.n353 2.13841
R9672 a_n13990_8177.n366 a_n13990_8177.n324 2.13841
R9673 a_n13990_8177.n231 a_n13990_8177.n178 2.0852
R9674 a_n13990_8177.n472 a_n13990_8177.n455 2.0852
R9675 a_n13990_8177.n556 a_n13990_8177.n304 1.95191
R9676 a_n13990_8177.n293 a_n13990_8177.n59 1.90397
R9677 a_n13990_8177.n557 a_n13990_8177.n556 1.80854
R9678 a_n13990_8177.n543 a_n13990_8177.n59 1.80603
R9679 a_n13990_8177.n355 a_n13990_8177.n333 1.73904
R9680 a_n13990_8177.n417 a_n13990_8177.n406 1.73904
R9681 a_n13990_8177.n530 a_n13990_8177.n304 1.73609
R9682 a_n13990_8177.n487 a_n13990_8177.n486 1.73609
R9683 a_n13990_8177.n292 a_n13990_8177.n291 1.65018
R9684 a_n13990_8177.n188 a_n13990_8177.n182 1.65018
R9685 a_n13990_8177.n542 a_n13990_8177.n303 1.56167
R9686 a_n13990_8177.n129 a_n13990_8177.n0 1.65553
R9687 a_n13990_8177.n559 a_n13990_8177.n3 1.65553
R9688 a_n13990_8177.n123 a_n13990_8177.n122 1.5005
R9689 a_n13990_8177.n240 a_n13990_8177.n239 1.5005
R9690 a_n13990_8177.n242 a_n13990_8177.n241 1.5005
R9691 a_n13990_8177.n302 a_n13990_8177.n301 1.5005
R9692 a_n13990_8177.n231 a_n13990_8177.n230 1.5005
R9693 a_n13990_8177.n267 a_n13990_8177.n167 1.5005
R9694 a_n13990_8177.n418 a_n13990_8177.n417 1.5005
R9695 a_n13990_8177.n397 a_n13990_8177.n396 1.5005
R9696 a_n13990_8177.n371 a_n13990_8177.n310 1.5005
R9697 a_n13990_8177.n355 a_n13990_8177.n354 1.5005
R9698 a_n13990_8177.n545 a_n13990_8177.n544 1.5005
R9699 a_n13990_8177.n555 a_n13990_8177.n554 1.5005
R9700 a_n13990_8177.n383 a_n13990_8177.n382 1.5005
R9701 a_n13990_8177.n381 a_n13990_8177.n380 1.5005
R9702 a_n13990_8177.n516 a_n13990_8177.n515 1.5005
R9703 a_n13990_8177.n474 a_n13990_8177.n473 1.5005
R9704 a_n13990_8177.n496 a_n13990_8177.n419 1.5005
R9705 a_n13990_8177.n541 a_n13990_8177.n540 1.5005
R9706 a_n13990_8177.n472 a_n13990_8177.n471 1.5005
R9707 a_n13990_8177.n559 a_n13990_8177.n558 1.5005
R9708 a_n13990_8177.n141 a_n13990_8177.n140 1.5005
R9709 a_n13990_8177.n130 a_n13990_8177.n129 1.5005
R9710 a_n13990_8177.n97 a_n13990_8177.n64 1.5005
R9711 a_n13990_8177.n166 a_n13990_8177.n165 1.5005
R9712 a_n13990_8177.n562 a_n13990_8177.n561 1.5005
R9713 a_n13990_8177.n571 a_n13990_8177.t225 1.4705
R9714 a_n13990_8177.n571 a_n13990_8177.n570 1.4705
R9715 a_n13990_8177.n154 a_n13990_8177.t212 1.4705
R9716 a_n13990_8177.n154 a_n13990_8177.n153 1.4705
R9717 a_n13990_8177.n156 a_n13990_8177.t154 1.4705
R9718 a_n13990_8177.n156 a_n13990_8177.n155 1.4705
R9719 a_n13990_8177.n147 a_n13990_8177.t134 1.4705
R9720 a_n13990_8177.n147 a_n13990_8177.n146 1.4705
R9721 a_n13990_8177.n149 a_n13990_8177.t119 1.4705
R9722 a_n13990_8177.n149 a_n13990_8177.n148 1.4705
R9723 a_n13990_8177.n53 a_n13990_8177.t122 1.4705
R9724 a_n13990_8177.n53 a_n13990_8177.n52 1.4705
R9725 a_n13990_8177.n55 a_n13990_8177.t178 1.4705
R9726 a_n13990_8177.n55 a_n13990_8177.n54 1.4705
R9727 a_n13990_8177.n66 a_n13990_8177.t198 1.4705
R9728 a_n13990_8177.n66 a_n13990_8177.n65 1.4705
R9729 a_n13990_8177.n71 a_n13990_8177.t250 1.4705
R9730 a_n13990_8177.n71 a_n13990_8177.n70 1.4705
R9731 a_n13990_8177.n86 a_n13990_8177.t137 1.4705
R9732 a_n13990_8177.n86 a_n13990_8177.n85 1.4705
R9733 a_n13990_8177.n88 a_n13990_8177.t146 1.4705
R9734 a_n13990_8177.n88 a_n13990_8177.n87 1.4705
R9735 a_n13990_8177.n99 a_n13990_8177.t237 1.4705
R9736 a_n13990_8177.n99 a_n13990_8177.n98 1.4705
R9737 a_n13990_8177.n101 a_n13990_8177.t245 1.4705
R9738 a_n13990_8177.n101 a_n13990_8177.n100 1.4705
R9739 a_n13990_8177.n111 a_n13990_8177.t149 1.4705
R9740 a_n13990_8177.n111 a_n13990_8177.n110 1.4705
R9741 a_n13990_8177.n113 a_n13990_8177.t162 1.4705
R9742 a_n13990_8177.n113 a_n13990_8177.n112 1.4705
R9743 a_n13990_8177.n79 a_n13990_8177.t227 1.4705
R9744 a_n13990_8177.n79 a_n13990_8177.n78 1.4705
R9745 a_n13990_8177.n81 a_n13990_8177.t235 1.4705
R9746 a_n13990_8177.n81 a_n13990_8177.n80 1.4705
R9747 a_n13990_8177.n128 a_n13990_8177.t224 1.4705
R9748 a_n13990_8177.n128 a_n13990_8177.n127 1.4705
R9749 a_n13990_8177.n126 a_n13990_8177.t232 1.4705
R9750 a_n13990_8177.n126 a_n13990_8177.n125 1.4705
R9751 a_n13990_8177.n137 a_n13990_8177.t94 1.4705
R9752 a_n13990_8177.n137 a_n13990_8177.n136 1.4705
R9753 a_n13990_8177.n134 a_n13990_8177.t147 1.4705
R9754 a_n13990_8177.n134 a_n13990_8177.n133 1.4705
R9755 a_n13990_8177.n63 a_n13990_8177.t249 1.4705
R9756 a_n13990_8177.n63 a_n13990_8177.n62 1.4705
R9757 a_n13990_8177.n61 a_n13990_8177.t190 1.4705
R9758 a_n13990_8177.n61 a_n13990_8177.n60 1.4705
R9759 a_n13990_8177.n177 a_n13990_8177.t37 1.4705
R9760 a_n13990_8177.n177 a_n13990_8177.n176 1.4705
R9761 a_n13990_8177.n181 a_n13990_8177.t70 1.4705
R9762 a_n13990_8177.n181 a_n13990_8177.n180 1.4705
R9763 a_n13990_8177.n245 a_n13990_8177.t311 1.4705
R9764 a_n13990_8177.n245 a_n13990_8177.n244 1.4705
R9765 a_n13990_8177.n247 a_n13990_8177.t310 1.4705
R9766 a_n13990_8177.n247 a_n13990_8177.n246 1.4705
R9767 a_n13990_8177.n250 a_n13990_8177.t48 1.4705
R9768 a_n13990_8177.n250 a_n13990_8177.n249 1.4705
R9769 a_n13990_8177.n252 a_n13990_8177.t330 1.4705
R9770 a_n13990_8177.n252 a_n13990_8177.n251 1.4705
R9771 a_n13990_8177.n256 a_n13990_8177.t329 1.4705
R9772 a_n13990_8177.n256 a_n13990_8177.n255 1.4705
R9773 a_n13990_8177.n258 a_n13990_8177.t328 1.4705
R9774 a_n13990_8177.n258 a_n13990_8177.n257 1.4705
R9775 a_n13990_8177.n262 a_n13990_8177.t12 1.4705
R9776 a_n13990_8177.n262 a_n13990_8177.n261 1.4705
R9777 a_n13990_8177.n264 a_n13990_8177.t21 1.4705
R9778 a_n13990_8177.n264 a_n13990_8177.n263 1.4705
R9779 a_n13990_8177.n269 a_n13990_8177.t15 1.4705
R9780 a_n13990_8177.n269 a_n13990_8177.n268 1.4705
R9781 a_n13990_8177.n271 a_n13990_8177.t13 1.4705
R9782 a_n13990_8177.n271 a_n13990_8177.n270 1.4705
R9783 a_n13990_8177.n275 a_n13990_8177.t35 1.4705
R9784 a_n13990_8177.n275 a_n13990_8177.n274 1.4705
R9785 a_n13990_8177.n277 a_n13990_8177.t34 1.4705
R9786 a_n13990_8177.n277 a_n13990_8177.n276 1.4705
R9787 a_n13990_8177.n281 a_n13990_8177.t8 1.4705
R9788 a_n13990_8177.n281 a_n13990_8177.n280 1.4705
R9789 a_n13990_8177.n283 a_n13990_8177.t7 1.4705
R9790 a_n13990_8177.n283 a_n13990_8177.n282 1.4705
R9791 a_n13990_8177.n287 a_n13990_8177.t30 1.4705
R9792 a_n13990_8177.n287 a_n13990_8177.n286 1.4705
R9793 a_n13990_8177.n289 a_n13990_8177.t29 1.4705
R9794 a_n13990_8177.n289 a_n13990_8177.n288 1.4705
R9795 a_n13990_8177.n208 a_n13990_8177.t51 1.4705
R9796 a_n13990_8177.n208 a_n13990_8177.n207 1.4705
R9797 a_n13990_8177.n210 a_n13990_8177.t52 1.4705
R9798 a_n13990_8177.n210 a_n13990_8177.n209 1.4705
R9799 a_n13990_8177.n213 a_n13990_8177.t1 1.4705
R9800 a_n13990_8177.n213 a_n13990_8177.n212 1.4705
R9801 a_n13990_8177.n215 a_n13990_8177.t331 1.4705
R9802 a_n13990_8177.n215 a_n13990_8177.n214 1.4705
R9803 a_n13990_8177.n219 a_n13990_8177.t308 1.4705
R9804 a_n13990_8177.n219 a_n13990_8177.n218 1.4705
R9805 a_n13990_8177.n221 a_n13990_8177.t309 1.4705
R9806 a_n13990_8177.n221 a_n13990_8177.n220 1.4705
R9807 a_n13990_8177.n225 a_n13990_8177.t313 1.4705
R9808 a_n13990_8177.n225 a_n13990_8177.n224 1.4705
R9809 a_n13990_8177.n227 a_n13990_8177.t314 1.4705
R9810 a_n13990_8177.n227 a_n13990_8177.n226 1.4705
R9811 a_n13990_8177.n202 a_n13990_8177.t49 1.4705
R9812 a_n13990_8177.n202 a_n13990_8177.n201 1.4705
R9813 a_n13990_8177.n204 a_n13990_8177.t50 1.4705
R9814 a_n13990_8177.n204 a_n13990_8177.n203 1.4705
R9815 a_n13990_8177.n196 a_n13990_8177.t9 1.4705
R9816 a_n13990_8177.n196 a_n13990_8177.n195 1.4705
R9817 a_n13990_8177.n198 a_n13990_8177.t11 1.4705
R9818 a_n13990_8177.n198 a_n13990_8177.n197 1.4705
R9819 a_n13990_8177.n190 a_n13990_8177.t347 1.4705
R9820 a_n13990_8177.n190 a_n13990_8177.n189 1.4705
R9821 a_n13990_8177.n192 a_n13990_8177.t349 1.4705
R9822 a_n13990_8177.n192 a_n13990_8177.n191 1.4705
R9823 a_n13990_8177.n184 a_n13990_8177.t14 1.4705
R9824 a_n13990_8177.n184 a_n13990_8177.n183 1.4705
R9825 a_n13990_8177.n186 a_n13990_8177.t16 1.4705
R9826 a_n13990_8177.n186 a_n13990_8177.n185 1.4705
R9827 a_n13990_8177.n299 a_n13990_8177.t45 1.4705
R9828 a_n13990_8177.n299 a_n13990_8177.n298 1.4705
R9829 a_n13990_8177.n295 a_n13990_8177.t351 1.4705
R9830 a_n13990_8177.n295 a_n13990_8177.n294 1.4705
R9831 a_n13990_8177.n174 a_n13990_8177.t43 1.4705
R9832 a_n13990_8177.n174 a_n13990_8177.n173 1.4705
R9833 a_n13990_8177.n171 a_n13990_8177.t336 1.4705
R9834 a_n13990_8177.n171 a_n13990_8177.n170 1.4705
R9835 a_n13990_8177.n237 a_n13990_8177.t350 1.4705
R9836 a_n13990_8177.n237 a_n13990_8177.n236 1.4705
R9837 a_n13990_8177.n233 a_n13990_8177.t312 1.4705
R9838 a_n13990_8177.n233 a_n13990_8177.n232 1.4705
R9839 a_n13990_8177.n553 a_n13990_8177.t136 1.4705
R9840 a_n13990_8177.n553 a_n13990_8177.n552 1.4705
R9841 a_n13990_8177.n550 a_n13990_8177.t108 1.4705
R9842 a_n13990_8177.n550 a_n13990_8177.n549 1.4705
R9843 a_n13990_8177.n547 a_n13990_8177.t248 1.4705
R9844 a_n13990_8177.n547 a_n13990_8177.n546 1.4705
R9845 a_n13990_8177.n308 a_n13990_8177.t159 1.4705
R9846 a_n13990_8177.n308 a_n13990_8177.n307 1.4705
R9847 a_n13990_8177.n322 a_n13990_8177.t155 1.4705
R9848 a_n13990_8177.n322 a_n13990_8177.n321 1.4705
R9849 a_n13990_8177.n345 a_n13990_8177.t255 1.4705
R9850 a_n13990_8177.n345 a_n13990_8177.n344 1.4705
R9851 a_n13990_8177.n351 a_n13990_8177.t167 1.4705
R9852 a_n13990_8177.n351 a_n13990_8177.n350 1.4705
R9853 a_n13990_8177.n336 a_n13990_8177.t239 1.4705
R9854 a_n13990_8177.n336 a_n13990_8177.n335 1.4705
R9855 a_n13990_8177.n361 a_n13990_8177.t182 1.4705
R9856 a_n13990_8177.n361 a_n13990_8177.n360 1.4705
R9857 a_n13990_8177.n363 a_n13990_8177.t194 1.4705
R9858 a_n13990_8177.n363 a_n13990_8177.n362 1.4705
R9859 a_n13990_8177.n329 a_n13990_8177.t233 1.4705
R9860 a_n13990_8177.n329 a_n13990_8177.n328 1.4705
R9861 a_n13990_8177.n331 a_n13990_8177.t240 1.4705
R9862 a_n13990_8177.n331 a_n13990_8177.n330 1.4705
R9863 a_n13990_8177.n379 a_n13990_8177.t177 1.4705
R9864 a_n13990_8177.n379 a_n13990_8177.n378 1.4705
R9865 a_n13990_8177.n376 a_n13990_8177.t105 1.4705
R9866 a_n13990_8177.n376 a_n13990_8177.n375 1.4705
R9867 a_n13990_8177.n373 a_n13990_8177.t189 1.4705
R9868 a_n13990_8177.n373 a_n13990_8177.n372 1.4705
R9869 a_n13990_8177.n369 a_n13990_8177.t265 1.4705
R9870 a_n13990_8177.n369 a_n13990_8177.n368 1.4705
R9871 a_n13990_8177.n319 a_n13990_8177.t226 1.4705
R9872 a_n13990_8177.n319 a_n13990_8177.n318 1.4705
R9873 a_n13990_8177.n388 a_n13990_8177.t152 1.4705
R9874 a_n13990_8177.n388 a_n13990_8177.n387 1.4705
R9875 a_n13990_8177.n394 a_n13990_8177.t236 1.4705
R9876 a_n13990_8177.n394 a_n13990_8177.n393 1.4705
R9877 a_n13990_8177.n313 a_n13990_8177.t139 1.4705
R9878 a_n13990_8177.n313 a_n13990_8177.n312 1.4705
R9879 a_n13990_8177.n408 a_n13990_8177.t251 1.4705
R9880 a_n13990_8177.n408 a_n13990_8177.n407 1.4705
R9881 a_n13990_8177.n410 a_n13990_8177.t142 1.4705
R9882 a_n13990_8177.n410 a_n13990_8177.n409 1.4705
R9883 a_n13990_8177.n402 a_n13990_8177.t130 1.4705
R9884 a_n13990_8177.n402 a_n13990_8177.n401 1.4705
R9885 a_n13990_8177.n404 a_n13990_8177.t215 1.4705
R9886 a_n13990_8177.n404 a_n13990_8177.n403 1.4705
R9887 a_n13990_8177.n466 a_n13990_8177.t302 1.4705
R9888 a_n13990_8177.n466 a_n13990_8177.n465 1.4705
R9889 a_n13990_8177.n468 a_n13990_8177.t303 1.4705
R9890 a_n13990_8177.n468 a_n13990_8177.n467 1.4705
R9891 a_n13990_8177.n457 a_n13990_8177.t321 1.4705
R9892 a_n13990_8177.n457 a_n13990_8177.n456 1.4705
R9893 a_n13990_8177.n459 a_n13990_8177.t323 1.4705
R9894 a_n13990_8177.n459 a_n13990_8177.n458 1.4705
R9895 a_n13990_8177.n529 a_n13990_8177.t320 1.4705
R9896 a_n13990_8177.n529 a_n13990_8177.n528 1.4705
R9897 a_n13990_8177.n532 a_n13990_8177.t345 1.4705
R9898 a_n13990_8177.n532 a_n13990_8177.n531 1.4705
R9899 a_n13990_8177.n535 a_n13990_8177.t90 1.4705
R9900 a_n13990_8177.n535 a_n13990_8177.n534 1.4705
R9901 a_n13990_8177.n538 a_n13990_8177.t58 1.4705
R9902 a_n13990_8177.n538 a_n13990_8177.n537 1.4705
R9903 a_n13990_8177.n526 a_n13990_8177.t59 1.4705
R9904 a_n13990_8177.n526 a_n13990_8177.n525 1.4705
R9905 a_n13990_8177.n523 a_n13990_8177.t283 1.4705
R9906 a_n13990_8177.n523 a_n13990_8177.n522 1.4705
R9907 a_n13990_8177.n520 a_n13990_8177.t80 1.4705
R9908 a_n13990_8177.n520 a_n13990_8177.n519 1.4705
R9909 a_n13990_8177.n518 a_n13990_8177.t82 1.4705
R9910 a_n13990_8177.n518 a_n13990_8177.n517 1.4705
R9911 a_n13990_8177.n504 a_n13990_8177.t91 1.4705
R9912 a_n13990_8177.n504 a_n13990_8177.n503 1.4705
R9913 a_n13990_8177.n502 a_n13990_8177.t298 1.4705
R9914 a_n13990_8177.n502 a_n13990_8177.n501 1.4705
R9915 a_n13990_8177.n500 a_n13990_8177.t269 1.4705
R9916 a_n13990_8177.n500 a_n13990_8177.n499 1.4705
R9917 a_n13990_8177.n498 a_n13990_8177.t322 1.4705
R9918 a_n13990_8177.n498 a_n13990_8177.n497 1.4705
R9919 a_n13990_8177.n495 a_n13990_8177.t318 1.4705
R9920 a_n13990_8177.n495 a_n13990_8177.n494 1.4705
R9921 a_n13990_8177.n493 a_n13990_8177.t54 1.4705
R9922 a_n13990_8177.n493 a_n13990_8177.n492 1.4705
R9923 a_n13990_8177.n491 a_n13990_8177.t273 1.4705
R9924 a_n13990_8177.n491 a_n13990_8177.n490 1.4705
R9925 a_n13990_8177.n489 a_n13990_8177.t280 1.4705
R9926 a_n13990_8177.n489 a_n13990_8177.n488 1.4705
R9927 a_n13990_8177.n485 a_n13990_8177.t285 1.4705
R9928 a_n13990_8177.n485 a_n13990_8177.n484 1.4705
R9929 a_n13990_8177.n482 a_n13990_8177.t276 1.4705
R9930 a_n13990_8177.n482 a_n13990_8177.n481 1.4705
R9931 a_n13990_8177.n479 a_n13990_8177.t85 1.4705
R9932 a_n13990_8177.n479 a_n13990_8177.n478 1.4705
R9933 a_n13990_8177.n476 a_n13990_8177.t292 1.4705
R9934 a_n13990_8177.n476 a_n13990_8177.n475 1.4705
R9935 a_n13990_8177.n437 a_n13990_8177.t278 1.4705
R9936 a_n13990_8177.n437 a_n13990_8177.n436 1.4705
R9937 a_n13990_8177.n434 a_n13990_8177.t268 1.4705
R9938 a_n13990_8177.n434 a_n13990_8177.n433 1.4705
R9939 a_n13990_8177.n431 a_n13990_8177.t317 1.4705
R9940 a_n13990_8177.n431 a_n13990_8177.n430 1.4705
R9941 a_n13990_8177.n429 a_n13990_8177.t53 1.4705
R9942 a_n13990_8177.n429 a_n13990_8177.n428 1.4705
R9943 a_n13990_8177.n454 a_n13990_8177.t0 1.4705
R9944 a_n13990_8177.n454 a_n13990_8177.n453 1.4705
R9945 a_n13990_8177.n452 a_n13990_8177.t343 1.4705
R9946 a_n13990_8177.n452 a_n13990_8177.n451 1.4705
R9947 a_n13990_8177.n450 a_n13990_8177.t299 1.4705
R9948 a_n13990_8177.n450 a_n13990_8177.n449 1.4705
R9949 a_n13990_8177.n448 a_n13990_8177.t324 1.4705
R9950 a_n13990_8177.n448 a_n13990_8177.n447 1.4705
R9951 a_n13990_8177.n446 a_n13990_8177.t55 1.4705
R9952 a_n13990_8177.n446 a_n13990_8177.n445 1.4705
R9953 a_n13990_8177.n444 a_n13990_8177.t81 1.4705
R9954 a_n13990_8177.n444 a_n13990_8177.n443 1.4705
R9955 a_n13990_8177.n442 a_n13990_8177.t301 1.4705
R9956 a_n13990_8177.n442 a_n13990_8177.n441 1.4705
R9957 a_n13990_8177.n440 a_n13990_8177.t60 1.4705
R9958 a_n13990_8177.n440 a_n13990_8177.n439 1.4705
R9959 a_n13990_8177.n510 a_n13990_8177.t339 1.4705
R9960 a_n13990_8177.n510 a_n13990_8177.n509 1.4705
R9961 a_n13990_8177.n512 a_n13990_8177.t338 1.4705
R9962 a_n13990_8177.n512 a_n13990_8177.n511 1.4705
R9963 a_n13990_8177.n421 a_n13990_8177.t83 1.4705
R9964 a_n13990_8177.n421 a_n13990_8177.n420 1.4705
R9965 a_n13990_8177.n423 a_n13990_8177.t319 1.4705
R9966 a_n13990_8177.n423 a_n13990_8177.n422 1.4705
R9967 a_n13990_8177.t267 a_n13990_8177.n573 1.4705
R9968 a_n13990_8177.n573 a_n13990_8177.n46 1.4705
R9969 a_n13990_8177.n158 a_n13990_8177.n157 1.46537
R9970 a_n13990_8177.n162 a_n13990_8177.n161 1.46537
R9971 a_n13990_8177.n151 a_n13990_8177.n150 1.46537
R9972 a_n13990_8177.n145 a_n13990_8177.n144 1.46537
R9973 a_n13990_8177.n48 a_n13990_8177.n47 1.46537
R9974 a_n13990_8177.n572 a_n13990_8177.n569 1.46537
R9975 a_n13990_8177.n568 a_n13990_8177.n567 1.46537
R9976 a_n13990_8177.n57 a_n13990_8177.n56 1.46537
R9977 a_n13990_8177.n90 a_n13990_8177.n89 1.46537
R9978 a_n13990_8177.n94 a_n13990_8177.n93 1.46537
R9979 a_n13990_8177.n103 a_n13990_8177.n102 1.46537
R9980 a_n13990_8177.n107 a_n13990_8177.n106 1.46537
R9981 a_n13990_8177.n109 a_n13990_8177.n108 1.46537
R9982 a_n13990_8177.n115 a_n13990_8177.n114 1.46537
R9983 a_n13990_8177.n119 a_n13990_8177.n118 1.46537
R9984 a_n13990_8177.n83 a_n13990_8177.n82 1.46537
R9985 a_n13990_8177.n365 a_n13990_8177.n364 1.46537
R9986 a_n13990_8177.n359 a_n13990_8177.n358 1.46537
R9987 a_n13990_8177.n333 a_n13990_8177.n332 1.46537
R9988 a_n13990_8177.n412 a_n13990_8177.n411 1.46537
R9989 a_n13990_8177.n416 a_n13990_8177.n415 1.46537
R9990 a_n13990_8177.n406 a_n13990_8177.n405 1.46537
R9991 a_n13990_8177.n464 a_n13990_8177.n463 1.46537
R9992 a_n13990_8177.n470 a_n13990_8177.n469 1.46537
R9993 a_n13990_8177.n462 a_n13990_8177.n461 1.46537
R9994 a_n13990_8177.n508 a_n13990_8177.n507 1.46537
R9995 a_n13990_8177.n514 a_n13990_8177.n513 1.46537
R9996 a_n13990_8177.n426 a_n13990_8177.n425 1.46537
R9997 a_n13990_8177.n254 a_n13990_8177.n253 1.46537
R9998 a_n13990_8177.n260 a_n13990_8177.n259 1.46537
R9999 a_n13990_8177.n266 a_n13990_8177.n265 1.46537
R10000 a_n13990_8177.n273 a_n13990_8177.n272 1.46537
R10001 a_n13990_8177.n279 a_n13990_8177.n278 1.46537
R10002 a_n13990_8177.n285 a_n13990_8177.n284 1.46537
R10003 a_n13990_8177.n291 a_n13990_8177.n290 1.46537
R10004 a_n13990_8177.n217 a_n13990_8177.n216 1.46537
R10005 a_n13990_8177.n223 a_n13990_8177.n222 1.46537
R10006 a_n13990_8177.n229 a_n13990_8177.n228 1.46537
R10007 a_n13990_8177.n206 a_n13990_8177.n205 1.46537
R10008 a_n13990_8177.n200 a_n13990_8177.n199 1.46537
R10009 a_n13990_8177.n194 a_n13990_8177.n193 1.46537
R10010 a_n13990_8177.n188 a_n13990_8177.n187 1.46537
R10011 a_n13990_8177.n164 a_n13990_8177.n163 1.46535
R10012 a_n13990_8177.n564 a_n13990_8177.n563 1.46535
R10013 a_n13990_8177.n96 a_n13990_8177.n95 1.46535
R10014 a_n13990_8177.n121 a_n13990_8177.n120 1.46535
R10015 a_n13990_8177.n542 a_n13990_8177.n541 1.34705
R10016 a_n13990_8177.n303 a_n13990_8177.n302 1.2981
R10017 a_n13990_8177.n558 a_n13990_8177.n557 1.27763
R10018 a_n13990_8177.n569 a_n13990_8177.n48 1.27228
R10019 a_n13990_8177.n74 a_n13990_8177.n72 1.27228
R10020 a_n13990_8177.n119 a_n13990_8177.n115 1.27228
R10021 a_n13990_8177.n115 a_n13990_8177.n109 1.27228
R10022 a_n13990_8177.n107 a_n13990_8177.n103 1.27228
R10023 a_n13990_8177.n94 a_n13990_8177.n90 1.27228
R10024 a_n13990_8177.n135 a_n13990_8177.n132 1.27228
R10025 a_n13990_8177.n352 a_n13990_8177.n349 1.27228
R10026 a_n13990_8177.n348 a_n13990_8177.n346 1.27228
R10027 a_n13990_8177.n365 a_n13990_8177.n359 1.27228
R10028 a_n13990_8177.n395 a_n13990_8177.n392 1.27228
R10029 a_n13990_8177.n391 a_n13990_8177.n389 1.27228
R10030 a_n13990_8177.n416 a_n13990_8177.n412 1.27228
R10031 a_n13990_8177.n569 a_n13990_8177.n568 1.27228
R10032 a_n13990_8177.n151 a_n13990_8177.n145 1.27228
R10033 a_n13990_8177.n162 a_n13990_8177.n158 1.27228
R10034 a_n13990_8177.n291 a_n13990_8177.n285 1.27228
R10035 a_n13990_8177.n279 a_n13990_8177.n273 1.27228
R10036 a_n13990_8177.n266 a_n13990_8177.n260 1.27228
R10037 a_n13990_8177.n194 a_n13990_8177.n188 1.27228
R10038 a_n13990_8177.n206 a_n13990_8177.n200 1.27228
R10039 a_n13990_8177.n229 a_n13990_8177.n223 1.27228
R10040 a_n13990_8177.n297 a_n13990_8177.n296 1.27228
R10041 a_n13990_8177.n235 a_n13990_8177.n234 1.27228
R10042 a_n13990_8177.n527 a_n13990_8177.n524 1.27228
R10043 a_n13990_8177.n539 a_n13990_8177.n536 1.27228
R10044 a_n13990_8177.n533 a_n13990_8177.n530 1.27228
R10045 a_n13990_8177.n438 a_n13990_8177.n435 1.27228
R10046 a_n13990_8177.n480 a_n13990_8177.n477 1.27228
R10047 a_n13990_8177.n486 a_n13990_8177.n483 1.27228
R10048 a_n13990_8177.n514 a_n13990_8177.n508 1.27228
R10049 a_n13990_8177.n470 a_n13990_8177.n464 1.27228
R10050 a_n13990_8177.n338 a_n13990_8177.n337 1.26756
R10051 a_n13990_8177.n346 a_n13990_8177.n343 1.26756
R10052 a_n13990_8177.n315 a_n13990_8177.n314 1.26756
R10053 a_n13990_8177.n389 a_n13990_8177.n386 1.26756
R10054 a_n13990_8177.n556 a_n13990_8177.n555 1.23567
R10055 a_n13990_8177.n544 a_n13990_8177.n543 1.23455
R10056 a_n13990_8177.n560 a_n13990_8177.n59 1.18682
R10057 a_n13990_8177.n69 a_n13990_8177.n68 1.01873
R10058 a_n13990_8177.n140 a_n13990_8177.n139 1.01873
R10059 a_n13990_8177.n473 a_n13990_8177.n419 0.822966
R10060 a_n13990_8177.n505 a_n13990_8177.n487 0.822966
R10061 a_n13990_8177.n353 a_n13990_8177.n340 0.796291
R10062 a_n13990_8177.n342 a_n13990_8177.n324 0.796291
R10063 a_n13990_8177.n396 a_n13990_8177.n317 0.796291
R10064 a_n13990_8177.n385 a_n13990_8177.n383 0.796291
R10065 a_n13990_8177.n354 a_n13990_8177.n310 0.780703
R10066 a_n13990_8177.n544 a_n13990_8177.n418 0.780703
R10067 a_n13990_8177.n381 a_n13990_8177.n366 0.780703
R10068 a_n13990_8177.n555 a_n13990_8177.n305 0.780703
R10069 a_n13990_8177.n124 a_n13990_8177.n123 0.778574
R10070 a_n13990_8177.n561 a_n13990_8177.n560 0.778574
R10071 a_n13990_8177.n130 a_n13990_8177.n64 0.778574
R10072 a_n13990_8177.n558 a_n13990_8177.n166 0.778574
R10073 a_n13990_8177.n561 a_n13990_8177.n58 0.738439
R10074 a_n13990_8177.n166 a_n13990_8177.n141 0.738439
R10075 a_n13990_8177.n293 a_n13990_8177.n292 0.737223
R10076 a_n13990_8177.n182 a_n13990_8177.n168 0.737223
R10077 a_n13990_8177.n302 a_n13990_8177.n167 0.737223
R10078 a_n13990_8177.n240 a_n13990_8177.n231 0.737223
R10079 a_n13990_8177.n243 a_n13990_8177.n168 0.725061
R10080 a_n13990_8177.n241 a_n13990_8177.n240 0.725061
R10081 a_n13990_8177.n122 a_n13990_8177.n121 0.699581
R10082 a_n13990_8177.n97 a_n13990_8177.n96 0.699581
R10083 a_n13990_8177.n564 a_n13990_8177.n562 0.699581
R10084 a_n13990_8177.n165 a_n13990_8177.n164 0.699581
R10085 a_n13990_8177.n541 a_n13990_8177.n516 0.639318
R10086 a_n13990_8177.n473 a_n13990_8177.n472 0.639318
R10087 a_n13990_8177.n506 a_n13990_8177.n304 0.639318
R10088 a_n13990_8177.n487 a_n13990_8177.n427 0.639318
R10089 a_n13990_8177.n418 a_n13990_8177.n397 0.638405
R10090 a_n13990_8177.n382 a_n13990_8177.n305 0.638405
R10091 a_n13990_8177.n397 a_n13990_8177.n310 0.628372
R10092 a_n13990_8177.n382 a_n13990_8177.n381 0.628372
R10093 a_n13990_8177.n543 a_n13990_8177.n542 0.606869
R10094 a_n13990_8177.n557 a_n13990_8177.n303 0.60536
R10095 a_n13990_8177.n292 a_n13990_8177.n243 0.585196
R10096 a_n13990_8177.n241 a_n13990_8177.n167 0.585196
R10097 a_n13990_8177.n516 a_n13990_8177.n419 0.585196
R10098 a_n13990_8177.n506 a_n13990_8177.n505 0.585196
R10099 a_n13990_8177.n122 a_n13990_8177.n83 0.557791
R10100 a_n13990_8177.n103 a_n13990_8177.n97 0.557791
R10101 a_n13990_8177.n562 a_n13990_8177.n57 0.557791
R10102 a_n13990_8177.n165 a_n13990_8177.n151 0.557791
R10103 a_n13990_8177.n124 a_n13990_8177.n58 0.530466
R10104 a_n13990_8177.n141 a_n13990_8177.n130 0.530466
R10105 a_n13990_8177.n353 a_n13990_8177.n352 0.476484
R10106 a_n13990_8177.n324 a_n13990_8177.n323 0.476484
R10107 a_n13990_8177.n396 a_n13990_8177.n395 0.476484
R10108 a_n13990_8177.n383 a_n13990_8177.n320 0.476484
R10109 a_n13990_8177.n28 a_n13990_8177.n371 0.478684
R10110 a_n13990_8177.n380 a_n13990_8177.n22 0.478684
R10111 a_n13990_8177.n18 a_n13990_8177.n545 0.478684
R10112 a_n13990_8177.n554 a_n13990_8177.n12 0.478684
R10113 a_n13990_8177.n540 a_n13990_8177.n527 0.236091
R10114 a_n13990_8177.n474 a_n13990_8177.n438 0.236091
R10115 a_n13990_8177.n267 a_n13990_8177.n266 0.150184
R10116 a_n13990_8177.n230 a_n13990_8177.n229 0.150184
R10117 a_n13990_8177.n1 a_n13990_8177.n2 1.27228
R10118 a_n13990_8177.n129 a_n13990_8177.n1 7.30549
R10119 a_n13990_8177.t103 a_n13990_8177.n0 6.96214
R10120 a_n13990_8177.n4 a_n13990_8177.n5 1.27228
R10121 a_n13990_8177.n559 a_n13990_8177.n4 7.30549
R10122 a_n13990_8177.t254 a_n13990_8177.n3 6.96214
R10123 a_n13990_8177.n10 a_n13990_8177.n11 1.26457
R10124 a_n13990_8177.n242 a_n13990_8177.n10 6.59229
R10125 a_n13990_8177.n174 a_n13990_8177.n9 5.10549
R10126 a_n13990_8177.n7 a_n13990_8177.n8 1.26457
R10127 a_n13990_8177.n178 a_n13990_8177.n7 6.59229
R10128 a_n13990_8177.n177 a_n13990_8177.n6 5.10549
R10129 a_n13990_8177.n30 a_n13990_8177.n31 1.27228
R10130 a_n13990_8177.n29 a_n13990_8177.n30 2.51878
R10131 a_n13990_8177.n371 a_n13990_8177.n29 0.794091
R10132 a_n13990_8177.n27 a_n13990_8177.n28 1.27228
R10133 a_n13990_8177.n26 a_n13990_8177.n27 2.60203
R10134 a_n13990_8177.n25 a_n13990_8177.n26 1.27228
R10135 a_n13990_8177.n24 a_n13990_8177.n25 1.27228
R10136 a_n13990_8177.n23 a_n13990_8177.n24 2.51878
R10137 a_n13990_8177.n380 a_n13990_8177.n23 0.794091
R10138 a_n13990_8177.t112 a_n13990_8177.n22 6.77266
R10139 a_n13990_8177.n20 a_n13990_8177.n21 1.27228
R10140 a_n13990_8177.n19 a_n13990_8177.n20 2.51878
R10141 a_n13990_8177.n545 a_n13990_8177.n19 0.794091
R10142 a_n13990_8177.n17 a_n13990_8177.n18 1.27228
R10143 a_n13990_8177.n16 a_n13990_8177.n17 2.60203
R10144 a_n13990_8177.n15 a_n13990_8177.n16 1.27228
R10145 a_n13990_8177.n14 a_n13990_8177.n15 1.27228
R10146 a_n13990_8177.n13 a_n13990_8177.n14 2.51878
R10147 a_n13990_8177.n554 a_n13990_8177.n13 0.794091
R10148 a_n13990_8177.t100 a_n13990_8177.n12 6.77266
R10149 a_n13990_8177.n37 a_n13990_8177.n38 3.79678
R10150 a_n13990_8177.n36 a_n13990_8177.n37 1.27228
R10151 a_n13990_8177.n496 a_n13990_8177.n36 0.238291
R10152 a_n13990_8177.n34 a_n13990_8177.n35 1.27228
R10153 a_n13990_8177.n33 a_n13990_8177.n34 3.79678
R10154 a_n13990_8177.n32 a_n13990_8177.n33 1.27228
R10155 a_n13990_8177.n505 a_n13990_8177.n32 1.73829
R10156 a_n13990_8177.n44 a_n13990_8177.n45 3.79678
R10157 a_n13990_8177.n43 a_n13990_8177.n44 1.27228
R10158 a_n13990_8177.n455 a_n13990_8177.n43 0.238291
R10159 a_n13990_8177.n41 a_n13990_8177.n42 1.27228
R10160 a_n13990_8177.n40 a_n13990_8177.n41 3.79678
R10161 a_n13990_8177.n39 a_n13990_8177.n40 1.27228
R10162 a_n13990_8177.n427 a_n13990_8177.n39 2.32299
R10163 a_n11317_n20927.t1 a_n11317_n20927.t7 23.2164
R10164 a_n11317_n20927.t5 a_n11317_n20927.t1 17.4491
R10165 a_n11317_n20927.t1 a_n11317_n20927.t4 17.1874
R10166 a_n11317_n20927.n0 a_n11317_n20927.t1 16.5634
R10167 VP.n11 VP.t25 8.38704
R10168 VP.n311 VP.t69 8.38704
R10169 VP.n125 VP.t7 8.37857
R10170 VP.n248 VP.t19 8.37857
R10171 VP.n58 VP.t60 8.31301
R10172 VP.n209 VP.t85 8.31301
R10173 VP.n388 VP.t5 8.29322
R10174 VP.n147 VP.t84 8.29322
R10175 VP.n387 VP.t3 8.10567
R10176 VP.n385 VP.t62 8.10567
R10177 VP.n384 VP.t81 8.10567
R10178 VP.n0 VP.t18 8.10567
R10179 VP.n339 VP.t47 8.10567
R10180 VP.n340 VP.t43 8.10567
R10181 VP.n322 VP.t40 8.10567
R10182 VP.n316 VP.t41 8.10567
R10183 VP.n310 VP.t13 8.10567
R10184 VP.n326 VP.t78 8.10567
R10185 VP.n325 VP.t20 8.10567
R10186 VP.n324 VP.t38 8.10567
R10187 VP.n332 VP.t65 8.10567
R10188 VP.n331 VP.t87 8.10567
R10189 VP.n369 VP.t54 8.10567
R10190 VP.n375 VP.t74 8.10567
R10191 VP.n116 VP.t46 8.10567
R10192 VP.n109 VP.t23 8.10567
R10193 VP.n103 VP.t4 8.10567
R10194 VP.n97 VP.t67 8.10567
R10195 VP.n120 VP.t30 8.10567
R10196 VP.n119 VP.t2 8.10567
R10197 VP.n118 VP.t32 8.10567
R10198 VP.n124 VP.t35 8.10567
R10199 VP.n123 VP.t76 8.10567
R10200 VP.n135 VP.t83 8.10567
R10201 VP.n53 VP.t11 8.10567
R10202 VP.n62 VP.t73 8.10567
R10203 VP.n57 VP.t66 8.10567
R10204 VP.n75 VP.t82 8.10567
R10205 VP.n74 VP.t55 8.10567
R10206 VP.n73 VP.t61 8.10567
R10207 VP.n95 VP.t64 8.10567
R10208 VP.n88 VP.t68 8.10567
R10209 VP.n81 VP.t22 8.10567
R10210 VP.n52 VP.t28 8.10567
R10211 VP.n39 VP.t44 8.10567
R10212 VP.n37 VP.t10 8.10567
R10213 VP.n36 VP.t72 8.10567
R10214 VP.n180 VP.t37 8.10567
R10215 VP.n161 VP.t29 8.10567
R10216 VP.n162 VP.t0 8.10567
R10217 VP.n163 VP.t31 8.10567
R10218 VP.n146 VP.t24 8.10567
R10219 VP.n144 VP.t12 8.10567
R10220 VP.n143 VP.t48 8.10567
R10221 VP.n22 VP.t71 8.10567
R10222 VP.n16 VP.t14 8.10567
R10223 VP.n10 VP.t51 8.10567
R10224 VP.n26 VP.t80 8.10567
R10225 VP.n25 VP.t53 8.10567
R10226 VP.n24 VP.t59 8.10567
R10227 VP.n32 VP.t27 8.10567
R10228 VP.n31 VP.t58 8.10567
R10229 VP.n192 VP.t50 8.10567
R10230 VP.n198 VP.t86 8.10567
R10231 VP.n242 VP.t34 8.10567
R10232 VP.n238 VP.t63 8.10567
R10233 VP.n237 VP.t26 8.10567
R10234 VP.n281 VP.t52 8.10567
R10235 VP.n261 VP.t16 8.10567
R10236 VP.n262 VP.t45 8.10567
R10237 VP.n263 VP.t42 8.10567
R10238 VP.n247 VP.t15 8.10567
R10239 VP.n245 VP.t75 8.10567
R10240 VP.n243 VP.t6 8.10567
R10241 VP.n223 VP.t56 8.10567
R10242 VP.n216 VP.t57 8.10567
R10243 VP.n210 VP.t33 8.10567
R10244 VP.n227 VP.t77 8.10567
R10245 VP.n226 VP.t17 8.10567
R10246 VP.n225 VP.t36 8.10567
R10247 VP.n283 VP.t79 8.10567
R10248 VP.n231 VP.t8 8.10567
R10249 VP.n230 VP.t70 8.10567
R10250 VP.n300 VP.t1 8.10567
R10251 VP.n342 VP.t21 8.10567
R10252 VP.n337 VP.t49 8.10567
R10253 VP.n336 VP.t9 8.10567
R10254 VP.n357 VP.t39 8.10567
R10255 VP.n381 VP.n380 7.37198
R10256 VP.n359 VP.n332 4.64261
R10257 VP.n182 VP.n32 4.64261
R10258 VP.n96 VP.n95 4.61892
R10259 VP.n284 VP.n283 4.61892
R10260 VP.n98 VP.n97 4.61655
R10261 VP.n282 VP.n281 4.61655
R10262 VP.n60 VP.n59 4.5005
R10263 VP.n61 VP.n56 4.5005
R10264 VP.n64 VP.n63 4.5005
R10265 VP.n65 VP.n55 4.5005
R10266 VP.n67 VP.n66 4.5005
R10267 VP.n68 VP.n54 4.5005
R10268 VP.n70 VP.n69 4.5005
R10269 VP.n72 VP.n71 4.5005
R10270 VP.n77 VP.n76 4.5005
R10271 VP.n79 VP.n78 4.5005
R10272 VP.n80 VP.n51 4.5005
R10273 VP.n83 VP.n82 4.5005
R10274 VP.n84 VP.n50 4.5005
R10275 VP.n86 VP.n85 4.5005
R10276 VP.n87 VP.n49 4.5005
R10277 VP.n90 VP.n89 4.5005
R10278 VP.n91 VP.n48 4.5005
R10279 VP.n93 VP.n92 4.5005
R10280 VP.n94 VP.n47 4.5005
R10281 VP.n99 VP.n46 4.5005
R10282 VP.n101 VP.n100 4.5005
R10283 VP.n102 VP.n45 4.5005
R10284 VP.n105 VP.n104 4.5005
R10285 VP.n106 VP.n44 4.5005
R10286 VP.n108 VP.n107 4.5005
R10287 VP.n110 VP.n43 4.5005
R10288 VP.n112 VP.n111 4.5005
R10289 VP.n113 VP.n42 4.5005
R10290 VP.n115 VP.n114 4.5005
R10291 VP.n117 VP.n40 4.5005
R10292 VP.n137 VP.n136 4.5005
R10293 VP.n134 VP.n41 4.5005
R10294 VP.n133 VP.n132 4.5005
R10295 VP.n131 VP.n121 4.5005
R10296 VP.n130 VP.n129 4.5005
R10297 VP.n128 VP.n122 4.5005
R10298 VP.n127 VP.n126 4.5005
R10299 VP.n23 VP.n5 4.5005
R10300 VP.n21 VP.n20 4.5005
R10301 VP.n19 VP.n7 4.5005
R10302 VP.n18 VP.n17 4.5005
R10303 VP.n15 VP.n8 4.5005
R10304 VP.n14 VP.n13 4.5005
R10305 VP.n12 VP.n9 4.5005
R10306 VP.n201 VP.n200 4.5005
R10307 VP.n199 VP.n6 4.5005
R10308 VP.n197 VP.n196 4.5005
R10309 VP.n195 VP.n27 4.5005
R10310 VP.n194 VP.n193 4.5005
R10311 VP.n191 VP.n28 4.5005
R10312 VP.n190 VP.n189 4.5005
R10313 VP.n188 VP.n29 4.5005
R10314 VP.n187 VP.n186 4.5005
R10315 VP.n185 VP.n30 4.5005
R10316 VP.n184 VP.n183 4.5005
R10317 VP.n165 VP.n164 4.5005
R10318 VP.n167 VP.n166 4.5005
R10319 VP.n168 VP.n38 4.5005
R10320 VP.n170 VP.n169 4.5005
R10321 VP.n172 VP.n171 4.5005
R10322 VP.n173 VP.n35 4.5005
R10323 VP.n175 VP.n174 4.5005
R10324 VP.n176 VP.n34 4.5005
R10325 VP.n178 VP.n177 4.5005
R10326 VP.n179 VP.n33 4.5005
R10327 VP.n160 VP.n159 4.5005
R10328 VP.n158 VP.n141 4.5005
R10329 VP.n157 VP.n156 4.5005
R10330 VP.n155 VP.n142 4.5005
R10331 VP.n154 VP.n153 4.5005
R10332 VP.n152 VP.n151 4.5005
R10333 VP.n150 VP.n145 4.5005
R10334 VP.n149 VP.n148 4.5005
R10335 VP.n212 VP.n211 4.5005
R10336 VP.n213 VP.n208 4.5005
R10337 VP.n215 VP.n214 4.5005
R10338 VP.n217 VP.n207 4.5005
R10339 VP.n219 VP.n218 4.5005
R10340 VP.n220 VP.n206 4.5005
R10341 VP.n222 VP.n221 4.5005
R10342 VP.n224 VP.n204 4.5005
R10343 VP.n302 VP.n301 4.5005
R10344 VP.n299 VP.n205 4.5005
R10345 VP.n298 VP.n297 4.5005
R10346 VP.n296 VP.n228 4.5005
R10347 VP.n295 VP.n294 4.5005
R10348 VP.n293 VP.n229 4.5005
R10349 VP.n292 VP.n291 4.5005
R10350 VP.n290 VP.n289 4.5005
R10351 VP.n288 VP.n232 4.5005
R10352 VP.n287 VP.n286 4.5005
R10353 VP.n285 VP.n233 4.5005
R10354 VP.n280 VP.n234 4.5005
R10355 VP.n279 VP.n278 4.5005
R10356 VP.n277 VP.n235 4.5005
R10357 VP.n276 VP.n275 4.5005
R10358 VP.n274 VP.n236 4.5005
R10359 VP.n273 VP.n272 4.5005
R10360 VP.n271 VP.n270 4.5005
R10361 VP.n269 VP.n239 4.5005
R10362 VP.n268 VP.n267 4.5005
R10363 VP.n266 VP.n240 4.5005
R10364 VP.n265 VP.n264 4.5005
R10365 VP.n260 VP.n259 4.5005
R10366 VP.n258 VP.n257 4.5005
R10367 VP.n256 VP.n244 4.5005
R10368 VP.n255 VP.n254 4.5005
R10369 VP.n253 VP.n252 4.5005
R10370 VP.n251 VP.n246 4.5005
R10371 VP.n250 VP.n249 4.5005
R10372 VP.n323 VP.n305 4.5005
R10373 VP.n321 VP.n320 4.5005
R10374 VP.n319 VP.n307 4.5005
R10375 VP.n318 VP.n317 4.5005
R10376 VP.n315 VP.n308 4.5005
R10377 VP.n314 VP.n313 4.5005
R10378 VP.n312 VP.n309 4.5005
R10379 VP.n378 VP.n377 4.5005
R10380 VP.n376 VP.n306 4.5005
R10381 VP.n374 VP.n373 4.5005
R10382 VP.n372 VP.n327 4.5005
R10383 VP.n371 VP.n370 4.5005
R10384 VP.n368 VP.n328 4.5005
R10385 VP.n367 VP.n366 4.5005
R10386 VP.n365 VP.n329 4.5005
R10387 VP.n364 VP.n363 4.5005
R10388 VP.n362 VP.n330 4.5005
R10389 VP.n361 VP.n360 4.5005
R10390 VP.n341 VP.n2 4.5005
R10391 VP.n344 VP.n343 4.5005
R10392 VP.n345 VP.n338 4.5005
R10393 VP.n347 VP.n346 4.5005
R10394 VP.n349 VP.n348 4.5005
R10395 VP.n350 VP.n335 4.5005
R10396 VP.n352 VP.n351 4.5005
R10397 VP.n353 VP.n334 4.5005
R10398 VP.n355 VP.n354 4.5005
R10399 VP.n356 VP.n333 4.5005
R10400 VP.n401 VP.n400 4.5005
R10401 VP.n399 VP.n1 4.5005
R10402 VP.n398 VP.n397 4.5005
R10403 VP.n396 VP.n383 4.5005
R10404 VP.n395 VP.n394 4.5005
R10405 VP.n393 VP.n392 4.5005
R10406 VP.n391 VP.n386 4.5005
R10407 VP.n390 VP.n389 4.5005
R10408 VP.n182 VP.n181 3.03856
R10409 VP.n359 VP.n358 3.03856
R10410 VP.n98 VP.n96 3.0245
R10411 VP.n284 VP.n282 3.0245
R10412 VP.n203 VP.n4 2.30989
R10413 VP.n139 VP.n138 2.30989
R10414 VP.n181 VP.n180 2.25752
R10415 VP.n358 VP.n357 2.25752
R10416 VP.n71 VP.n4 2.18975
R10417 VP.n138 VP.n40 2.18975
R10418 VP.n303 VP.n204 2.18975
R10419 VP.n265 VP.n241 2.18975
R10420 VP.n202 VP.n5 2.16725
R10421 VP.n165 VP.n140 2.16725
R10422 VP.n379 VP.n305 2.16725
R10423 VP.n382 VP.n2 2.16725
R10424 VP.n304 VP.n303 1.5005
R10425 VP.n203 VP.n202 1.5005
R10426 VP.n241 VP.n3 1.5005
R10427 VP.n140 VP.n139 1.5005
R10428 VP.n382 VP.n381 1.5005
R10429 VP.n380 VP.n379 1.5005
R10430 VP.n148 VP.n147 1.392
R10431 VP.n389 VP.n388 1.392
R10432 VP.n59 VP.n58 1.38741
R10433 VP.n212 VP.n209 1.38741
R10434 VP.n136 VP.n120 1.24866
R10435 VP.n76 VP.n75 1.24866
R10436 VP.n261 VP.n260 1.24866
R10437 VP.n301 VP.n227 1.24866
R10438 VP.n118 VP.n117 1.24629
R10439 VP.n73 VP.n72 1.24629
R10440 VP.n264 VP.n263 1.24629
R10441 VP.n225 VP.n224 1.24629
R10442 VP.n304 VP.n203 1.23709
R10443 VP.n139 VP.n3 1.23709
R10444 VP.n324 VP.n323 1.22261
R10445 VP.n164 VP.n163 1.22261
R10446 VP.n24 VP.n23 1.22261
R10447 VP.n341 VP.n340 1.22261
R10448 VP.n377 VP.n326 1.21313
R10449 VP.n161 VP.n160 1.21313
R10450 VP.n200 VP.n26 1.21313
R10451 VP.n12 VP.n11 1.12904
R10452 VP.n312 VP.n311 1.12904
R10453 VP.n126 VP.n125 1.11862
R10454 VP.n249 VP.n248 1.11862
R10455 VP VP.n0 1.06037
R10456 VP.n380 VP.n304 0.809892
R10457 VP.n381 VP.n3 0.809892
R10458 VP.n77 VP.n4 0.752
R10459 VP.n138 VP.n137 0.752
R10460 VP.n303 VP.n302 0.752
R10461 VP.n259 VP.n241 0.752
R10462 VP.n202 VP.n201 0.71825
R10463 VP.n159 VP.n140 0.71825
R10464 VP.n379 VP.n378 0.71825
R10465 VP.n400 VP.n382 0.71825
R10466 VP.n325 VP.n324 0.673132
R10467 VP.n326 VP.n325 0.673132
R10468 VP.n119 VP.n118 0.673132
R10469 VP.n120 VP.n119 0.673132
R10470 VP.n74 VP.n73 0.673132
R10471 VP.n75 VP.n74 0.673132
R10472 VP.n163 VP.n162 0.673132
R10473 VP.n162 VP.n161 0.673132
R10474 VP.n25 VP.n24 0.673132
R10475 VP.n26 VP.n25 0.673132
R10476 VP.n263 VP.n262 0.673132
R10477 VP.n262 VP.n261 0.673132
R10478 VP.n226 VP.n225 0.673132
R10479 VP.n227 VP.n226 0.673132
R10480 VP.n340 VP.n339 0.673132
R10481 VP.n339 VP.n0 0.673132
R10482 VP.n147 VP.n146 0.45279
R10483 VP.n388 VP.n387 0.45279
R10484 VP.n58 VP.n57 0.430924
R10485 VP.n210 VP.n209 0.430924
R10486 VP.n128 VP.n127 0.394842
R10487 VP.n108 VP.n44 0.394842
R10488 VP.n87 VP.n86 0.394842
R10489 VP.n63 VP.n61 0.394842
R10490 VP.n251 VP.n250 0.394842
R10491 VP.n274 VP.n273 0.394842
R10492 VP.n293 VP.n292 0.394842
R10493 VP.n215 VP.n208 0.394842
R10494 VP.n133 VP.n121 0.381816
R10495 VP.n102 VP.n101 0.381816
R10496 VP.n82 VP.n80 0.381816
R10497 VP.n256 VP.n255 0.381816
R10498 VP.n279 VP.n235 0.381816
R10499 VP.n298 VP.n228 0.381816
R10500 VP.n374 VP.n327 0.379447
R10501 VP.n368 VP.n367 0.379447
R10502 VP.n363 VP.n362 0.379447
R10503 VP.n314 VP.n309 0.379447
R10504 VP.n317 VP.n307 0.379447
R10505 VP.n156 VP.n155 0.379447
R10506 VP.n151 VP.n150 0.379447
R10507 VP.n179 VP.n178 0.379447
R10508 VP.n174 VP.n173 0.379447
R10509 VP.n169 VP.n168 0.379447
R10510 VP.n197 VP.n27 0.379447
R10511 VP.n191 VP.n190 0.379447
R10512 VP.n186 VP.n185 0.379447
R10513 VP.n14 VP.n9 0.379447
R10514 VP.n17 VP.n7 0.379447
R10515 VP.n356 VP.n355 0.379447
R10516 VP.n351 VP.n350 0.379447
R10517 VP.n346 VP.n345 0.379447
R10518 VP.n397 VP.n396 0.379447
R10519 VP.n392 VP.n391 0.379447
R10520 VP.n64 VP.n56 0.375125
R10521 VP.n85 VP.n49 0.375125
R10522 VP.n107 VP.n106 0.375125
R10523 VP.n126 VP.n122 0.375125
R10524 VP.n214 VP.n213 0.375125
R10525 VP.n291 VP.n229 0.375125
R10526 VP.n272 VP.n236 0.375125
R10527 VP.n249 VP.n246 0.375125
R10528 VP.n83 VP.n51 0.36275
R10529 VP.n100 VP.n45 0.36275
R10530 VP.n132 VP.n131 0.36275
R10531 VP.n297 VP.n296 0.36275
R10532 VP.n278 VP.n277 0.36275
R10533 VP.n254 VP.n244 0.36275
R10534 VP.n13 VP.n12 0.3605
R10535 VP.n19 VP.n18 0.3605
R10536 VP.n196 VP.n195 0.3605
R10537 VP.n189 VP.n28 0.3605
R10538 VP.n187 VP.n30 0.3605
R10539 VP.n177 VP.n33 0.3605
R10540 VP.n175 VP.n35 0.3605
R10541 VP.n170 VP.n38 0.3605
R10542 VP.n157 VP.n142 0.3605
R10543 VP.n152 VP.n145 0.3605
R10544 VP.n313 VP.n312 0.3605
R10545 VP.n319 VP.n318 0.3605
R10546 VP.n373 VP.n372 0.3605
R10547 VP.n366 VP.n328 0.3605
R10548 VP.n364 VP.n330 0.3605
R10549 VP.n354 VP.n333 0.3605
R10550 VP.n352 VP.n335 0.3605
R10551 VP.n347 VP.n338 0.3605
R10552 VP.n398 VP.n383 0.3605
R10553 VP.n393 VP.n386 0.3605
R10554 VP.n125 VP.n124 0.348488
R10555 VP.n248 VP.n247 0.348488
R10556 VP.n311 VP.n310 0.327481
R10557 VP.n11 VP.n10 0.327481
R10558 VP.n111 VP.n42 0.302474
R10559 VP.n93 VP.n48 0.302474
R10560 VP.n68 VP.n67 0.302474
R10561 VP.n269 VP.n268 0.302474
R10562 VP.n288 VP.n287 0.302474
R10563 VP.n218 VP.n206 0.302474
R10564 VP.n66 VP.n54 0.287375
R10565 VP.n92 VP.n91 0.287375
R10566 VP.n113 VP.n112 0.287375
R10567 VP.n220 VP.n219 0.287375
R10568 VP.n286 VP.n232 0.287375
R10569 VP.n267 VP.n239 0.287375
R10570 VP.n181 VP.n33 0.208099
R10571 VP.n358 VP.n333 0.208099
R10572 VP VP.n401 0.153263
R10573 VP.n377 VP.n376 0.147342
R10574 VP.n370 VP.n327 0.147342
R10575 VP.n367 VP.n329 0.147342
R10576 VP.n362 VP.n361 0.147342
R10577 VP.n315 VP.n314 0.147342
R10578 VP.n321 VP.n307 0.147342
R10579 VP.n134 VP.n133 0.147342
R10580 VP.n129 VP.n128 0.147342
R10581 VP.n101 VP.n46 0.147342
R10582 VP.n104 VP.n44 0.147342
R10583 VP.n111 VP.n110 0.147342
R10584 VP.n115 VP.n42 0.147342
R10585 VP.n80 VP.n79 0.147342
R10586 VP.n86 VP.n50 0.147342
R10587 VP.n89 VP.n48 0.147342
R10588 VP.n94 VP.n93 0.147342
R10589 VP.n61 VP.n60 0.147342
R10590 VP.n67 VP.n55 0.147342
R10591 VP.n69 VP.n68 0.147342
R10592 VP.n160 VP.n141 0.147342
R10593 VP.n155 VP.n154 0.147342
R10594 VP.n150 VP.n149 0.147342
R10595 VP.n178 VP.n34 0.147342
R10596 VP.n173 VP.n172 0.147342
R10597 VP.n168 VP.n167 0.147342
R10598 VP.n200 VP.n199 0.147342
R10599 VP.n193 VP.n27 0.147342
R10600 VP.n190 VP.n29 0.147342
R10601 VP.n185 VP.n184 0.147342
R10602 VP.n15 VP.n14 0.147342
R10603 VP.n21 VP.n7 0.147342
R10604 VP.n257 VP.n256 0.147342
R10605 VP.n252 VP.n251 0.147342
R10606 VP.n280 VP.n279 0.147342
R10607 VP.n275 VP.n274 0.147342
R10608 VP.n270 VP.n269 0.147342
R10609 VP.n268 VP.n240 0.147342
R10610 VP.n299 VP.n298 0.147342
R10611 VP.n294 VP.n293 0.147342
R10612 VP.n289 VP.n288 0.147342
R10613 VP.n287 VP.n233 0.147342
R10614 VP.n211 VP.n208 0.147342
R10615 VP.n218 VP.n217 0.147342
R10616 VP.n222 VP.n206 0.147342
R10617 VP.n355 VP.n334 0.147342
R10618 VP.n350 VP.n349 0.147342
R10619 VP.n345 VP.n344 0.147342
R10620 VP.n401 VP.n1 0.147342
R10621 VP.n396 VP.n395 0.147342
R10622 VP.n391 VP.n390 0.147342
R10623 VP.n375 VP.n374 0.142605
R10624 VP.n369 VP.n368 0.142605
R10625 VP.n363 VP.n331 0.142605
R10626 VP.n310 VP.n309 0.142605
R10627 VP.n317 VP.n316 0.142605
R10628 VP.n323 VP.n322 0.142605
R10629 VP.n156 VP.n143 0.142605
R10630 VP.n151 VP.n144 0.142605
R10631 VP.n180 VP.n179 0.142605
R10632 VP.n174 VP.n36 0.142605
R10633 VP.n169 VP.n37 0.142605
R10634 VP.n164 VP.n39 0.142605
R10635 VP.n198 VP.n197 0.142605
R10636 VP.n192 VP.n191 0.142605
R10637 VP.n186 VP.n31 0.142605
R10638 VP.n10 VP.n9 0.142605
R10639 VP.n17 VP.n16 0.142605
R10640 VP.n23 VP.n22 0.142605
R10641 VP.n357 VP.n356 0.142605
R10642 VP.n351 VP.n336 0.142605
R10643 VP.n346 VP.n337 0.142605
R10644 VP.n342 VP.n341 0.142605
R10645 VP.n397 VP.n384 0.142605
R10646 VP.n392 VP.n385 0.142605
R10647 VP.n59 VP.n56 0.14
R10648 VP.n65 VP.n64 0.14
R10649 VP.n66 VP.n65 0.14
R10650 VP.n70 VP.n54 0.14
R10651 VP.n71 VP.n70 0.14
R10652 VP.n78 VP.n77 0.14
R10653 VP.n78 VP.n51 0.14
R10654 VP.n84 VP.n83 0.14
R10655 VP.n85 VP.n84 0.14
R10656 VP.n90 VP.n49 0.14
R10657 VP.n91 VP.n90 0.14
R10658 VP.n92 VP.n47 0.14
R10659 VP.n96 VP.n47 0.14
R10660 VP.n99 VP.n98 0.14
R10661 VP.n100 VP.n99 0.14
R10662 VP.n105 VP.n45 0.14
R10663 VP.n106 VP.n105 0.14
R10664 VP.n107 VP.n43 0.14
R10665 VP.n112 VP.n43 0.14
R10666 VP.n114 VP.n113 0.14
R10667 VP.n114 VP.n40 0.14
R10668 VP.n137 VP.n41 0.14
R10669 VP.n132 VP.n41 0.14
R10670 VP.n131 VP.n130 0.14
R10671 VP.n130 VP.n122 0.14
R10672 VP.n13 VP.n8 0.14
R10673 VP.n18 VP.n8 0.14
R10674 VP.n20 VP.n19 0.14
R10675 VP.n20 VP.n5 0.14
R10676 VP.n201 VP.n6 0.14
R10677 VP.n196 VP.n6 0.14
R10678 VP.n195 VP.n194 0.14
R10679 VP.n194 VP.n28 0.14
R10680 VP.n189 VP.n188 0.14
R10681 VP.n188 VP.n187 0.14
R10682 VP.n183 VP.n30 0.14
R10683 VP.n183 VP.n182 0.14
R10684 VP.n177 VP.n176 0.14
R10685 VP.n176 VP.n175 0.14
R10686 VP.n171 VP.n35 0.14
R10687 VP.n171 VP.n170 0.14
R10688 VP.n166 VP.n38 0.14
R10689 VP.n166 VP.n165 0.14
R10690 VP.n159 VP.n158 0.14
R10691 VP.n158 VP.n157 0.14
R10692 VP.n153 VP.n142 0.14
R10693 VP.n153 VP.n152 0.14
R10694 VP.n148 VP.n145 0.14
R10695 VP.n213 VP.n212 0.14
R10696 VP.n214 VP.n207 0.14
R10697 VP.n219 VP.n207 0.14
R10698 VP.n221 VP.n220 0.14
R10699 VP.n221 VP.n204 0.14
R10700 VP.n302 VP.n205 0.14
R10701 VP.n297 VP.n205 0.14
R10702 VP.n296 VP.n295 0.14
R10703 VP.n295 VP.n229 0.14
R10704 VP.n291 VP.n290 0.14
R10705 VP.n290 VP.n232 0.14
R10706 VP.n286 VP.n285 0.14
R10707 VP.n285 VP.n284 0.14
R10708 VP.n282 VP.n234 0.14
R10709 VP.n278 VP.n234 0.14
R10710 VP.n277 VP.n276 0.14
R10711 VP.n276 VP.n236 0.14
R10712 VP.n272 VP.n271 0.14
R10713 VP.n271 VP.n239 0.14
R10714 VP.n267 VP.n266 0.14
R10715 VP.n266 VP.n265 0.14
R10716 VP.n259 VP.n258 0.14
R10717 VP.n258 VP.n244 0.14
R10718 VP.n254 VP.n253 0.14
R10719 VP.n253 VP.n246 0.14
R10720 VP.n313 VP.n308 0.14
R10721 VP.n318 VP.n308 0.14
R10722 VP.n320 VP.n319 0.14
R10723 VP.n320 VP.n305 0.14
R10724 VP.n378 VP.n306 0.14
R10725 VP.n373 VP.n306 0.14
R10726 VP.n372 VP.n371 0.14
R10727 VP.n371 VP.n328 0.14
R10728 VP.n366 VP.n365 0.14
R10729 VP.n365 VP.n364 0.14
R10730 VP.n360 VP.n330 0.14
R10731 VP.n360 VP.n359 0.14
R10732 VP.n354 VP.n353 0.14
R10733 VP.n353 VP.n352 0.14
R10734 VP.n348 VP.n335 0.14
R10735 VP.n348 VP.n347 0.14
R10736 VP.n343 VP.n338 0.14
R10737 VP.n343 VP.n2 0.14
R10738 VP.n400 VP.n399 0.14
R10739 VP.n399 VP.n398 0.14
R10740 VP.n394 VP.n383 0.14
R10741 VP.n394 VP.n393 0.14
R10742 VP.n389 VP.n386 0.14
R10743 VP.n117 VP.n116 0.118921
R10744 VP.n72 VP.n53 0.118921
R10745 VP.n264 VP.n242 0.118921
R10746 VP.n224 VP.n223 0.118921
R10747 VP.n136 VP.n135 0.116553
R10748 VP.n76 VP.n52 0.116553
R10749 VP.n260 VP.n243 0.116553
R10750 VP.n301 VP.n300 0.116553
R10751 VP.n123 VP.n121 0.114184
R10752 VP.n103 VP.n102 0.114184
R10753 VP.n82 VP.n81 0.114184
R10754 VP.n255 VP.n245 0.114184
R10755 VP.n237 VP.n235 0.114184
R10756 VP.n230 VP.n228 0.114184
R10757 VP.n127 VP.n124 0.0987895
R10758 VP.n109 VP.n108 0.0987895
R10759 VP.n88 VP.n87 0.0987895
R10760 VP.n63 VP.n62 0.0987895
R10761 VP.n250 VP.n247 0.0987895
R10762 VP.n273 VP.n238 0.0987895
R10763 VP.n292 VP.n231 0.0987895
R10764 VP.n216 VP.n215 0.0987895
R10765 VP.n110 VP.n109 0.0490526
R10766 VP.n89 VP.n88 0.0490526
R10767 VP.n62 VP.n55 0.0490526
R10768 VP.n270 VP.n238 0.0490526
R10769 VP.n289 VP.n231 0.0490526
R10770 VP.n217 VP.n216 0.0490526
R10771 VP.n129 VP.n123 0.0336579
R10772 VP.n104 VP.n103 0.0336579
R10773 VP.n81 VP.n50 0.0336579
R10774 VP.n60 VP.n57 0.0336579
R10775 VP.n252 VP.n245 0.0336579
R10776 VP.n275 VP.n237 0.0336579
R10777 VP.n294 VP.n230 0.0336579
R10778 VP.n211 VP.n210 0.0336579
R10779 VP.n135 VP.n134 0.0312895
R10780 VP.n97 VP.n46 0.0312895
R10781 VP.n79 VP.n52 0.0312895
R10782 VP.n257 VP.n243 0.0312895
R10783 VP.n281 VP.n280 0.0312895
R10784 VP.n300 VP.n299 0.0312895
R10785 VP.n116 VP.n115 0.0289211
R10786 VP.n95 VP.n94 0.0289211
R10787 VP.n69 VP.n53 0.0289211
R10788 VP.n242 VP.n240 0.0289211
R10789 VP.n283 VP.n233 0.0289211
R10790 VP.n223 VP.n222 0.0289211
R10791 VP.n376 VP.n375 0.00523684
R10792 VP.n370 VP.n369 0.00523684
R10793 VP.n331 VP.n329 0.00523684
R10794 VP.n361 VP.n332 0.00523684
R10795 VP.n316 VP.n315 0.00523684
R10796 VP.n322 VP.n321 0.00523684
R10797 VP.n143 VP.n141 0.00523684
R10798 VP.n154 VP.n144 0.00523684
R10799 VP.n149 VP.n146 0.00523684
R10800 VP.n36 VP.n34 0.00523684
R10801 VP.n172 VP.n37 0.00523684
R10802 VP.n167 VP.n39 0.00523684
R10803 VP.n199 VP.n198 0.00523684
R10804 VP.n193 VP.n192 0.00523684
R10805 VP.n31 VP.n29 0.00523684
R10806 VP.n184 VP.n32 0.00523684
R10807 VP.n16 VP.n15 0.00523684
R10808 VP.n22 VP.n21 0.00523684
R10809 VP.n336 VP.n334 0.00523684
R10810 VP.n349 VP.n337 0.00523684
R10811 VP.n344 VP.n342 0.00523684
R10812 VP.n384 VP.n1 0.00523684
R10813 VP.n395 VP.n385 0.00523684
R10814 VP.n390 VP.n387 0.00523684
R10815 a_n13990_n6451.n202 a_n13990_n6451.n201 8.18538
R10816 a_n13990_n6451.n83 a_n13990_n6451.n79 7.22198
R10817 a_n13990_n6451.n229 a_n13990_n6451.n228 7.22198
R10818 a_n13990_n6451.n61 a_n13990_n6451.n58 6.77653
R10819 a_n13990_n6451.n29 a_n13990_n6451.n26 6.77653
R10820 a_n13990_n6451.n117 a_n13990_n6451.t122 6.7761
R10821 a_n13990_n6451.n47 a_n13990_n6451.t134 6.7761
R10822 a_n13990_n6451.n25 a_n13990_n6451.n133 6.86989
R10823 a_n13990_n6451.n9 a_n13990_n6451.n91 6.77231
R10824 a_n13990_n6451.n19 a_n13990_n6451.n203 6.77231
R10825 a_n13990_n6451.n196 a_n13990_n6451.n193 6.53862
R10826 a_n13990_n6451.n217 a_n13990_n6451.n202 5.95467
R10827 a_n13990_n6451.n152 a_n13990_n6451.n148 5.89898
R10828 a_n13990_n6451.n172 a_n13990_n6451.t20 5.66511
R10829 a_n13990_n6451.n162 a_n13990_n6451.t21 5.66511
R10830 a_n13990_n6451.n174 a_n13990_n6451.n173 5.66379
R10831 a_n13990_n6451.n164 a_n13990_n6451.n163 5.66379
R10832 a_n13990_n6451.n162 a_n13990_n6451.n161 5.65285
R10833 a_n13990_n6451.n143 a_n13990_n6451.n142 5.61877
R10834 a_n13990_n6451.n145 a_n13990_n6451.n144 5.61877
R10835 a_n13990_n6451.n137 a_n13990_n6451.n136 5.61877
R10836 a_n13990_n6451.n112 a_n13990_n6451.t107 5.50607
R10837 a_n13990_n6451.n30 a_n13990_n6451.t85 5.50607
R10838 a_n13990_n6451.n67 a_n13990_n6451.t95 5.50607
R10839 a_n13990_n6451.n62 a_n13990_n6451.t130 5.50607
R10840 a_n13990_n6451.n114 a_n13990_n6451.n113 5.50475
R10841 a_n13990_n6451.n108 a_n13990_n6451.n107 5.50475
R10842 a_n13990_n6451.n106 a_n13990_n6451.t62 5.50475
R10843 a_n13990_n6451.n66 a_n13990_n6451.n65 5.50475
R10844 a_n13990_n6451.n72 a_n13990_n6451.n71 5.50475
R10845 a_n13990_n6451.n73 a_n13990_n6451.t77 5.50475
R10846 a_n13990_n6451.n64 a_n13990_n6451.n63 5.50475
R10847 a_n13990_n6451.n234 a_n13990_n6451.n233 5.50475
R10848 a_n13990_n6451.n200 a_n13990_n6451.t26 5.28484
R10849 a_n13990_n6451.n22 a_n13990_n6451.n181 5.29079
R10850 a_n13990_n6451.n177 a_n13990_n6451.n176 4.88835
R10851 a_n13990_n6451.n123 a_n13990_n6451.n122 4.88517
R10852 a_n13990_n6451.n183 a_n13990_n6451.n21 4.02009
R10853 a_n13990_n6451.t36 a_n13990_n6451.n20 5.28011
R10854 a_n13990_n6451.t41 a_n13990_n6451.n22 5.28011
R10855 a_n13990_n6451.n0 a_n13990_n6451.n103 4.0312
R10856 a_n13990_n6451.n101 a_n13990_n6451.n1 5.5012
R10857 a_n13990_n6451.t97 a_n13990_n6451.n2 5.5012
R10858 a_n13990_n6451.n100 a_n13990_n6451.n3 4.0312
R10859 a_n13990_n6451.n98 a_n13990_n6451.n4 5.5012
R10860 a_n13990_n6451.t114 a_n13990_n6451.n5 5.5012
R10861 a_n13990_n6451.n97 a_n13990_n6451.n6 4.0312
R10862 a_n13990_n6451.n94 a_n13990_n6451.n7 5.5012
R10863 a_n13990_n6451.t70 a_n13990_n6451.n8 5.5012
R10864 a_n13990_n6451.n93 a_n13990_n6451.n9 4.0312
R10865 a_n13990_n6451.n10 a_n13990_n6451.n215 4.0312
R10866 a_n13990_n6451.n213 a_n13990_n6451.n11 5.5012
R10867 a_n13990_n6451.t120 a_n13990_n6451.n12 5.5012
R10868 a_n13990_n6451.n212 a_n13990_n6451.n13 4.0312
R10869 a_n13990_n6451.n210 a_n13990_n6451.n14 5.5012
R10870 a_n13990_n6451.t76 a_n13990_n6451.n15 5.5012
R10871 a_n13990_n6451.n209 a_n13990_n6451.n16 4.0312
R10872 a_n13990_n6451.n206 a_n13990_n6451.n17 5.5012
R10873 a_n13990_n6451.t101 a_n13990_n6451.n18 5.5012
R10874 a_n13990_n6451.n205 a_n13990_n6451.n19 4.0312
R10875 a_n13990_n6451.n23 a_n13990_n6451.n141 4.40099
R10876 a_n13990_n6451.n24 a_n13990_n6451.n139 4.40099
R10877 a_n13990_n6451.n135 a_n13990_n6451.n25 4.40099
R10878 a_n13990_n6451.n171 a_n13990_n6451.n170 4.40379
R10879 a_n13990_n6451.n168 a_n13990_n6451.n167 4.40379
R10880 a_n13990_n6451.n151 a_n13990_n6451.n150 4.40142
R10881 a_n13990_n6451.n126 a_n13990_n6451.n125 4.40142
R10882 a_n13990_n6451.n82 a_n13990_n6451.n81 4.24002
R10883 a_n13990_n6451.n51 a_n13990_n6451.n50 4.24002
R10884 a_n13990_n6451.n227 a_n13990_n6451.n226 4.24002
R10885 a_n13990_n6451.n38 a_n13990_n6451.n37 4.24002
R10886 a_n13990_n6451.n190 a_n13990_n6451.t39 4.22616
R10887 a_n13990_n6451.n117 a_n13990_n6451.n116 4.03475
R10888 a_n13990_n6451.n111 a_n13990_n6451.n110 4.03475
R10889 a_n13990_n6451.n33 a_n13990_n6451.n32 4.03475
R10890 a_n13990_n6451.n29 a_n13990_n6451.n28 4.03475
R10891 a_n13990_n6451.n47 a_n13990_n6451.n46 4.03475
R10892 a_n13990_n6451.n70 a_n13990_n6451.n69 4.03475
R10893 a_n13990_n6451.n76 a_n13990_n6451.n75 4.03475
R10894 a_n13990_n6451.n61 a_n13990_n6451.n60 4.03475
R10895 a_n13990_n6451.n199 a_n13990_n6451.n198 4.02484
R10896 a_n13990_n6451.n196 a_n13990_n6451.n195 4.02484
R10897 a_n13990_n6451.n190 a_n13990_n6451.t33 4.02247
R10898 a_n13990_n6451.n192 a_n13990_n6451.n191 3.96014
R10899 a_n13990_n6451.n179 a_n13990_n6451.n120 3.94195
R10900 a_n13990_n6451.n151 a_n13990_n6451.n149 3.84721
R10901 a_n13990_n6451.n126 a_n13990_n6451.n124 3.84721
R10902 a_n13990_n6451.n171 a_n13990_n6451.n168 3.81703
R10903 a_n13990_n6451.n199 a_n13990_n6451.n196 3.80578
R10904 a_n13990_n6451.n82 a_n13990_n6451.n80 3.68818
R10905 a_n13990_n6451.n51 a_n13990_n6451.n49 3.68818
R10906 a_n13990_n6451.n227 a_n13990_n6451.n225 3.68818
R10907 a_n13990_n6451.n38 a_n13990_n6451.n36 3.68818
R10908 a_n13990_n6451.n90 a_n13990_n6451.n89 3.23904
R10909 a_n13990_n6451.n224 a_n13990_n6451.n218 3.23904
R10910 a_n13990_n6451.n159 a_n13990_n6451.n158 3.23004
R10911 a_n13990_n6451.n157 a_n13990_n6451.n156 3.14142
R10912 a_n13990_n6451.n131 a_n13990_n6451.n130 3.14142
R10913 a_n13990_n6451.n189 a_n13990_n6451.n186 2.96616
R10914 a_n13990_n6451.n88 a_n13990_n6451.n87 2.77002
R10915 a_n13990_n6451.n56 a_n13990_n6451.n55 2.77002
R10916 a_n13990_n6451.n223 a_n13990_n6451.n222 2.77002
R10917 a_n13990_n6451.n43 a_n13990_n6451.n42 2.77002
R10918 a_n13990_n6451.n189 a_n13990_n6451.n188 2.76247
R10919 a_n13990_n6451.n57 a_n13990_n6451.n51 2.73714
R10920 a_n13990_n6451.n44 a_n13990_n6451.n38 2.73714
R10921 a_n13990_n6451.n191 a_n13990_n6451.n189 2.71914
R10922 a_n13990_n6451.n132 a_n13990_n6451.n126 2.71914
R10923 a_n13990_n6451.n179 a_n13990_n6451.n178 2.64424
R10924 a_n13990_n6451.n73 a_n13990_n6451.n72 2.60203
R10925 a_n13990_n6451.n108 a_n13990_n6451.n106 2.60203
R10926 a_n13990_n6451.n157 a_n13990_n6451.n154 2.58721
R10927 a_n13990_n6451.n131 a_n13990_n6451.n128 2.58721
R10928 a_n13990_n6451.n164 a_n13990_n6451.n162 2.55136
R10929 a_n13990_n6451.n174 a_n13990_n6451.n172 2.55136
R10930 a_n13990_n6451.n233 a_n13990_n6451.n30 2.52471
R10931 a_n13990_n6451.n64 a_n13990_n6451.n62 2.52436
R10932 a_n13990_n6451.n67 a_n13990_n6451.n66 2.52436
R10933 a_n13990_n6451.n114 a_n13990_n6451.n112 2.52436
R10934 a_n13990_n6451.n147 a_n13990_n6451.n146 2.2807
R10935 a_n13990_n6451.n159 a_n13990_n6451.n123 2.2807
R10936 a_n13990_n6451.n88 a_n13990_n6451.n85 2.21818
R10937 a_n13990_n6451.n56 a_n13990_n6451.n53 2.21818
R10938 a_n13990_n6451.n223 a_n13990_n6451.n220 2.21818
R10939 a_n13990_n6451.n43 a_n13990_n6451.n40 2.21818
R10940 a_n13990_n6451.n78 a_n13990_n6451.n77 2.13841
R10941 a_n13990_n6451.n90 a_n13990_n6451.n48 2.13841
R10942 a_n13990_n6451.n79 a_n13990_n6451.n57 1.73904
R10943 a_n13990_n6451.n229 a_n13990_n6451.n44 1.73904
R10944 a_n13990_n6451.n201 a_n13990_n6451.n200 1.73609
R10945 a_n13990_n6451.n148 a_n13990_n6451.n132 1.73004
R10946 a_n13990_n6451.n207 a_n13990_n6451.n35 1.5005
R10947 a_n13990_n6451.n230 a_n13990_n6451.n229 1.5005
R10948 a_n13990_n6451.n95 a_n13990_n6451.n34 1.5005
R10949 a_n13990_n6451.n79 a_n13990_n6451.n78 1.5005
R10950 a_n13990_n6451.n148 a_n13990_n6451.n147 1.5005
R10951 a_n13990_n6451.n165 a_n13990_n6451.n120 1.5005
R10952 a_n13990_n6451.n178 a_n13990_n6451.n177 1.5005
R10953 a_n13990_n6451.n217 a_n13990_n6451.n216 1.5005
R10954 a_n13990_n6451.n105 a_n13990_n6451.n104 1.5005
R10955 a_n13990_n6451.n119 a_n13990_n6451.n118 1.5005
R10956 a_n13990_n6451.n232 a_n13990_n6451.n231 1.5005
R10957 a_n13990_n6451.n116 a_n13990_n6451.t66 1.4705
R10958 a_n13990_n6451.n116 a_n13990_n6451.n115 1.4705
R10959 a_n13990_n6451.n110 a_n13990_n6451.t115 1.4705
R10960 a_n13990_n6451.n110 a_n13990_n6451.n109 1.4705
R10961 a_n13990_n6451.n32 a_n13990_n6451.t71 1.4705
R10962 a_n13990_n6451.n32 a_n13990_n6451.n31 1.4705
R10963 a_n13990_n6451.n28 a_n13990_n6451.t108 1.4705
R10964 a_n13990_n6451.n28 a_n13990_n6451.n27 1.4705
R10965 a_n13990_n6451.n46 a_n13990_n6451.t65 1.4705
R10966 a_n13990_n6451.n46 a_n13990_n6451.n45 1.4705
R10967 a_n13990_n6451.n69 a_n13990_n6451.t137 1.4705
R10968 a_n13990_n6451.n69 a_n13990_n6451.n68 1.4705
R10969 a_n13990_n6451.n75 a_n13990_n6451.t119 1.4705
R10970 a_n13990_n6451.n75 a_n13990_n6451.n74 1.4705
R10971 a_n13990_n6451.n60 a_n13990_n6451.t75 1.4705
R10972 a_n13990_n6451.n60 a_n13990_n6451.n59 1.4705
R10973 a_n13990_n6451.n85 a_n13990_n6451.t139 1.4705
R10974 a_n13990_n6451.n85 a_n13990_n6451.n84 1.4705
R10975 a_n13990_n6451.n87 a_n13990_n6451.t141 1.4705
R10976 a_n13990_n6451.n87 a_n13990_n6451.n86 1.4705
R10977 a_n13990_n6451.n53 a_n13990_n6451.t86 1.4705
R10978 a_n13990_n6451.n53 a_n13990_n6451.n52 1.4705
R10979 a_n13990_n6451.n55 a_n13990_n6451.t88 1.4705
R10980 a_n13990_n6451.n55 a_n13990_n6451.n54 1.4705
R10981 a_n13990_n6451.n103 a_n13990_n6451.t129 1.4705
R10982 a_n13990_n6451.n103 a_n13990_n6451.n102 1.4705
R10983 a_n13990_n6451.n100 a_n13990_n6451.t69 1.4705
R10984 a_n13990_n6451.n100 a_n13990_n6451.n99 1.4705
R10985 a_n13990_n6451.n97 a_n13990_n6451.t91 1.4705
R10986 a_n13990_n6451.n97 a_n13990_n6451.n96 1.4705
R10987 a_n13990_n6451.n93 a_n13990_n6451.t90 1.4705
R10988 a_n13990_n6451.n93 a_n13990_n6451.n92 1.4705
R10989 a_n13990_n6451.n220 a_n13990_n6451.t96 1.4705
R10990 a_n13990_n6451.n220 a_n13990_n6451.n219 1.4705
R10991 a_n13990_n6451.n222 a_n13990_n6451.t94 1.4705
R10992 a_n13990_n6451.n222 a_n13990_n6451.n221 1.4705
R10993 a_n13990_n6451.n40 a_n13990_n6451.t124 1.4705
R10994 a_n13990_n6451.n40 a_n13990_n6451.n39 1.4705
R10995 a_n13990_n6451.n42 a_n13990_n6451.t121 1.4705
R10996 a_n13990_n6451.n42 a_n13990_n6451.n41 1.4705
R10997 a_n13990_n6451.n215 a_n13990_n6451.t79 1.4705
R10998 a_n13990_n6451.n215 a_n13990_n6451.n214 1.4705
R10999 a_n13990_n6451.n212 a_n13990_n6451.t132 1.4705
R11000 a_n13990_n6451.n212 a_n13990_n6451.n211 1.4705
R11001 a_n13990_n6451.n209 a_n13990_n6451.t87 1.4705
R11002 a_n13990_n6451.n209 a_n13990_n6451.n208 1.4705
R11003 a_n13990_n6451.n205 a_n13990_n6451.t128 1.4705
R11004 a_n13990_n6451.n205 a_n13990_n6451.n204 1.4705
R11005 a_n13990_n6451.n89 a_n13990_n6451.n88 1.46537
R11006 a_n13990_n6451.n83 a_n13990_n6451.n82 1.46537
R11007 a_n13990_n6451.n57 a_n13990_n6451.n56 1.46537
R11008 a_n13990_n6451.n224 a_n13990_n6451.n223 1.46537
R11009 a_n13990_n6451.n228 a_n13990_n6451.n227 1.46537
R11010 a_n13990_n6451.n44 a_n13990_n6451.n43 1.46537
R11011 a_n13990_n6451.n158 a_n13990_n6451.n157 1.46537
R11012 a_n13990_n6451.n152 a_n13990_n6451.n151 1.46537
R11013 a_n13990_n6451.n132 a_n13990_n6451.n131 1.46537
R11014 a_n13990_n6451.n191 a_n13990_n6451.n190 1.46537
R11015 a_n13990_n6451.n202 a_n13990_n6451.n35 1.37875
R11016 a_n13990_n6451.n76 a_n13990_n6451.n73 1.27228
R11017 a_n13990_n6451.n72 a_n13990_n6451.n70 1.27228
R11018 a_n13990_n6451.n89 a_n13990_n6451.n83 1.27228
R11019 a_n13990_n6451.n228 a_n13990_n6451.n224 1.27228
R11020 a_n13990_n6451.n106 a_n13990_n6451.n33 1.27228
R11021 a_n13990_n6451.n111 a_n13990_n6451.n108 1.27228
R11022 a_n13990_n6451.n62 a_n13990_n6451.n61 1.26756
R11023 a_n13990_n6451.n70 a_n13990_n6451.n67 1.26756
R11024 a_n13990_n6451.n30 a_n13990_n6451.n29 1.26756
R11025 a_n13990_n6451.n112 a_n13990_n6451.n111 1.26756
R11026 a_n13990_n6451.n184 a_n13990_n6451.n179 1.26344
R11027 a_n13990_n6451.n198 a_n13990_n6451.t27 1.2605
R11028 a_n13990_n6451.n198 a_n13990_n6451.n197 1.2605
R11029 a_n13990_n6451.n195 a_n13990_n6451.t35 1.2605
R11030 a_n13990_n6451.n195 a_n13990_n6451.n194 1.2605
R11031 a_n13990_n6451.n183 a_n13990_n6451.t37 1.2605
R11032 a_n13990_n6451.n183 a_n13990_n6451.n182 1.2605
R11033 a_n13990_n6451.n181 a_n13990_n6451.t42 1.2605
R11034 a_n13990_n6451.n181 a_n13990_n6451.n180 1.2605
R11035 a_n13990_n6451.n186 a_n13990_n6451.t40 1.2605
R11036 a_n13990_n6451.n186 a_n13990_n6451.n185 1.2605
R11037 a_n13990_n6451.n188 a_n13990_n6451.t34 1.2605
R11038 a_n13990_n6451.n188 a_n13990_n6451.n187 1.2605
R11039 a_n13990_n6451.n122 a_n13990_n6451.t19 1.2605
R11040 a_n13990_n6451.n122 a_n13990_n6451.n121 1.2605
R11041 a_n13990_n6451.n141 a_n13990_n6451.t46 1.2605
R11042 a_n13990_n6451.n141 a_n13990_n6451.n140 1.2605
R11043 a_n13990_n6451.n139 a_n13990_n6451.t12 1.2605
R11044 a_n13990_n6451.n139 a_n13990_n6451.n138 1.2605
R11045 a_n13990_n6451.n135 a_n13990_n6451.t53 1.2605
R11046 a_n13990_n6451.n135 a_n13990_n6451.n134 1.2605
R11047 a_n13990_n6451.n176 a_n13990_n6451.t10 1.2605
R11048 a_n13990_n6451.n176 a_n13990_n6451.n175 1.2605
R11049 a_n13990_n6451.n170 a_n13990_n6451.t52 1.2605
R11050 a_n13990_n6451.n170 a_n13990_n6451.n169 1.2605
R11051 a_n13990_n6451.n167 a_n13990_n6451.t3 1.2605
R11052 a_n13990_n6451.n167 a_n13990_n6451.n166 1.2605
R11053 a_n13990_n6451.n161 a_n13990_n6451.t16 1.2605
R11054 a_n13990_n6451.n161 a_n13990_n6451.n160 1.2605
R11055 a_n13990_n6451.n154 a_n13990_n6451.t51 1.2605
R11056 a_n13990_n6451.n154 a_n13990_n6451.n153 1.2605
R11057 a_n13990_n6451.n156 a_n13990_n6451.t24 1.2605
R11058 a_n13990_n6451.n156 a_n13990_n6451.n155 1.2605
R11059 a_n13990_n6451.n128 a_n13990_n6451.t11 1.2605
R11060 a_n13990_n6451.n128 a_n13990_n6451.n127 1.2605
R11061 a_n13990_n6451.n130 a_n13990_n6451.t8 1.2605
R11062 a_n13990_n6451.n130 a_n13990_n6451.n129 1.2605
R11063 a_n13990_n6451.n158 a_n13990_n6451.n152 1.25428
R11064 a_n13990_n6451.n200 a_n13990_n6451.n199 1.25428
R11065 a_n13990_n6451.n172 a_n13990_n6451.n171 1.24956
R11066 a_n13990_n6451.n145 a_n13990_n6451.n23 1.25162
R11067 a_n13990_n6451.n77 a_n13990_n6451.n64 0.796291
R11068 a_n13990_n6451.n66 a_n13990_n6451.n48 0.796291
R11069 a_n13990_n6451.n118 a_n13990_n6451.n114 0.796291
R11070 a_n13990_n6451.n233 a_n13990_n6451.n232 0.795934
R11071 a_n13990_n6451.n78 a_n13990_n6451.n34 0.780703
R11072 a_n13990_n6451.n230 a_n13990_n6451.n35 0.780703
R11073 a_n13990_n6451.n105 a_n13990_n6451.n90 0.780703
R11074 a_n13990_n6451.n218 a_n13990_n6451.n217 0.780703
R11075 a_n13990_n6451.n165 a_n13990_n6451.n164 0.769291
R11076 a_n13990_n6451.n177 a_n13990_n6451.n174 0.769291
R11077 a_n13990_n6451.n146 a_n13990_n6451.n137 0.767125
R11078 a_n13990_n6451.n143 a_n13990_n6451.n123 0.767125
R11079 a_n13990_n6451.n201 a_n13990_n6451.n192 0.639318
R11080 a_n13990_n6451.n231 a_n13990_n6451.n230 0.638405
R11081 a_n13990_n6451.n147 a_n13990_n6451.n120 0.638405
R11082 a_n13990_n6451.n178 a_n13990_n6451.n159 0.638405
R11083 a_n13990_n6451.n218 a_n13990_n6451.n119 0.638405
R11084 a_n13990_n6451.n231 a_n13990_n6451.n34 0.628372
R11085 a_n13990_n6451.n119 a_n13990_n6451.n105 0.628372
R11086 a_n13990_n6451.n192 a_n13990_n6451.n184 0.585196
R11087 a_n13990_n6451.n168 a_n13990_n6451.n165 0.485484
R11088 a_n13990_n6451.n77 a_n13990_n6451.n76 0.476484
R11089 a_n13990_n6451.n48 a_n13990_n6451.n47 0.476484
R11090 a_n13990_n6451.n232 a_n13990_n6451.n33 0.476484
R11091 a_n13990_n6451.n118 a_n13990_n6451.n117 0.476484
R11092 a_n13990_n6451.n146 a_n13990_n6451.n24 0.484998
R11093 a_n13990_n6451.n6 a_n13990_n6451.n95 0.478684
R11094 a_n13990_n6451.n104 a_n13990_n6451.n0 0.478684
R11095 a_n13990_n6451.n16 a_n13990_n6451.n207 0.478684
R11096 a_n13990_n6451.n216 a_n13990_n6451.n10 0.478684
R11097 a_n13990_n6451.n8 a_n13990_n6451.n9 1.27228
R11098 a_n13990_n6451.n7 a_n13990_n6451.n8 2.51878
R11099 a_n13990_n6451.n95 a_n13990_n6451.n7 0.794091
R11100 a_n13990_n6451.n5 a_n13990_n6451.n6 1.27228
R11101 a_n13990_n6451.n4 a_n13990_n6451.n5 2.60203
R11102 a_n13990_n6451.n3 a_n13990_n6451.n4 1.27228
R11103 a_n13990_n6451.n2 a_n13990_n6451.n3 1.27228
R11104 a_n13990_n6451.n1 a_n13990_n6451.n2 2.51878
R11105 a_n13990_n6451.n104 a_n13990_n6451.n1 0.794091
R11106 a_n13990_n6451.t57 a_n13990_n6451.n0 6.77266
R11107 a_n13990_n6451.n18 a_n13990_n6451.n19 1.27228
R11108 a_n13990_n6451.n17 a_n13990_n6451.n18 2.51878
R11109 a_n13990_n6451.n207 a_n13990_n6451.n17 0.794091
R11110 a_n13990_n6451.n15 a_n13990_n6451.n16 1.27228
R11111 a_n13990_n6451.n14 a_n13990_n6451.n15 2.60203
R11112 a_n13990_n6451.n13 a_n13990_n6451.n14 1.27228
R11113 a_n13990_n6451.n12 a_n13990_n6451.n13 1.27228
R11114 a_n13990_n6451.n11 a_n13990_n6451.n12 2.51878
R11115 a_n13990_n6451.n216 a_n13990_n6451.n11 0.794091
R11116 a_n13990_n6451.t136 a_n13990_n6451.n10 6.77266
R11117 a_n13990_n6451.n21 a_n13990_n6451.n22 3.15817
R11118 a_n13990_n6451.n20 a_n13990_n6451.n21 1.27188
R11119 a_n13990_n6451.n184 a_n13990_n6451.n20 1.73829
R11120 a_n13990_n6451.n137 a_n13990_n6451.n25 3.17898
R11121 a_n13990_n6451.n145 a_n13990_n6451.n24 3.19023
R11122 a_n13990_n6451.n143 a_n13990_n6451.n23 3.17898
R11123 VN.n0 VN.t28 8.10567
R11124 VN.n754 VN.t45 8.10567
R11125 VN.n36 VN.t12 8.10567
R11126 VN.n30 VN.t6 8.10567
R11127 VN.n49 VN.t62 8.10567
R11128 VN.n55 VN.t1 8.10567
R11129 VN.n786 VN.t67 8.10567
R11130 VN.n779 VN.t4 8.10567
R11131 VN.n835 VN.t58 8.10567
R11132 VN.n841 VN.t81 8.10567
R11133 VN.n190 VN.t21 8.10567
R11134 VN.n349 VN.t14 8.10567
R11135 VN.n343 VN.t38 8.10567
R11136 VN.n338 VN.t85 8.10567
R11137 VN.n333 VN.t2 8.10567
R11138 VN.n316 VN.t54 8.10567
R11139 VN.n305 VN.t31 8.10567
R11140 VN.n296 VN.t11 8.10567
R11141 VN.n287 VN.t72 8.10567
R11142 VN.n172 VN.t66 8.10567
R11143 VN.n267 VN.t75 8.10567
R11144 VN.n180 VN.t29 8.10567
R11145 VN.n184 VN.t34 8.10567
R11146 VN.n330 VN.t18 8.10567
R11147 VN.n323 VN.t80 8.10567
R11148 VN.n156 VN.t19 8.10567
R11149 VN.n246 VN.t69 8.10567
R11150 VN.n239 VN.t42 8.10567
R11151 VN.n188 VN.t51 8.10567
R11152 VN.n194 VN.t78 8.10567
R11153 VN.n212 VN.t70 8.10567
R11154 VN.n202 VN.t60 8.10567
R11155 VN.n100 VN.t20 8.10567
R11156 VN.n404 VN.t13 8.10567
R11157 VN.n398 VN.t37 8.10567
R11158 VN.n393 VN.t83 8.10567
R11159 VN.n389 VN.t0 8.10567
R11160 VN.n381 VN.t52 8.10567
R11161 VN.n144 VN.t30 8.10567
R11162 VN.n451 VN.t7 8.10567
R11163 VN.n457 VN.t71 8.10567
R11164 VN.n133 VN.t63 8.10567
R11165 VN.n126 VN.t73 8.10567
R11166 VN.n121 VN.t27 8.10567
R11167 VN.n478 VN.t33 8.10567
R11168 VN.n387 VN.t48 8.10567
R11169 VN.n386 VN.t17 8.10567
R11170 VN.n436 VN.t43 8.10567
R11171 VN.n114 VN.t82 8.10567
R11172 VN.n107 VN.t46 8.10567
R11173 VN.n65 VN.t84 8.10567
R11174 VN.n72 VN.t77 8.10567
R11175 VN.n74 VN.t68 8.10567
R11176 VN.n78 VN.t59 8.10567
R11177 VN.n532 VN.t44 8.10567
R11178 VN.n606 VN.t9 8.10567
R11179 VN.n600 VN.t5 8.10567
R11180 VN.n595 VN.t61 8.10567
R11181 VN.n590 VN.t87 8.10567
R11182 VN.n650 VN.t26 8.10567
R11183 VN.n660 VN.t55 8.10567
R11184 VN.n669 VN.t15 8.10567
R11185 VN.n678 VN.t40 8.10567
R11186 VN.n566 VN.t65 8.10567
R11187 VN.n559 VN.t3 8.10567
R11188 VN.n554 VN.t57 8.10567
R11189 VN.n549 VN.t79 8.10567
R11190 VN.n586 VN.t24 8.10567
R11191 VN.n585 VN.t53 8.10567
R11192 VN.n646 VN.t50 8.10567
R11193 VN.n546 VN.t86 8.10567
R11194 VN.n539 VN.t25 8.10567
R11195 VN.n489 VN.t39 8.10567
R11196 VN.n521 VN.t47 8.10567
R11197 VN.n512 VN.t22 8.10567
R11198 VN.n503 VN.t74 8.10567
R11199 VN.n743 VN.t49 8.10567
R11200 VN.n727 VN.t23 8.10567
R11201 VN.n730 VN.t76 8.10567
R11202 VN.n19 VN.t8 8.10567
R11203 VN.n12 VN.t36 8.10567
R11204 VN.n7 VN.t35 8.10567
R11205 VN.n768 VN.t64 8.10567
R11206 VN.n761 VN.t10 8.10567
R11207 VN.n719 VN.t32 8.10567
R11208 VN.n798 VN.t56 8.10567
R11209 VN.n793 VN.t16 8.10567
R11210 VN.n819 VN.t41 8.10567
R11211 VN.n846 VN.n845 7.83574
R11212 VN.n204 VN.n201 4.65575
R11213 VN.n505 VN.n502 4.65575
R11214 VN.n350 VN.n345 4.64641
R11215 VN.n607 VN.n604 4.64641
R11216 VN.n351 VN.n350 4.64
R11217 VN.n79 VN.n77 4.64
R11218 VN.n406 VN.n405 4.64
R11219 VN.n80 VN.n79 4.64
R11220 VN.n407 VN.n406 4.64
R11221 VN.n610 VN.n604 4.64
R11222 VN.n733 VN.n732 4.64
R11223 VN.n38 VN.n37 4.64
R11224 VN.n732 VN.n731 4.64
R11225 VN.n39 VN.n38 4.64
R11226 VN.n426 VN.n387 4.54125
R11227 VN.n115 VN.n114 4.54125
R11228 VN.n20 VN.n19 4.54125
R11229 VN.n769 VN.n768 4.54125
R11230 VN.n331 VN.n330 4.53893
R11231 VN.n247 VN.n246 4.53893
R11232 VN.n636 VN.n586 4.53893
R11233 VN.n547 VN.n546 4.53893
R11234 VN.n377 VN.n376 4.51011
R11235 VN.n284 VN.n170 4.51011
R11236 VN.n250 VN.n248 4.51011
R11237 VN.n634 VN.n589 4.51011
R11238 VN.n681 VN.n680 4.51011
R11239 VN.n711 VN.n710 4.51011
R11240 VN.n317 VN.n150 4.50691
R11241 VN.n283 VN.n282 4.50691
R11242 VN.n233 VN.n232 4.50691
R11243 VN.n649 VN.n580 4.50691
R11244 VN.n683 VN.n682 4.50691
R11245 VN.n533 VN.n483 4.50691
R11246 VN.n245 VN.n185 4.5005
R11247 VN.n244 VN.n243 4.5005
R11248 VN.n242 VN.n186 4.5005
R11249 VN.n241 VN.n240 4.5005
R11250 VN.n238 VN.n187 4.5005
R11251 VN.n237 VN.n236 4.5005
R11252 VN.n329 VN.n153 4.5005
R11253 VN.n328 VN.n327 4.5005
R11254 VN.n326 VN.n154 4.5005
R11255 VN.n325 VN.n324 4.5005
R11256 VN.n322 VN.n155 4.5005
R11257 VN.n321 VN.n320 4.5005
R11258 VN.n251 VN.n250 4.5005
R11259 VN.n253 VN.n252 4.5005
R11260 VN.n182 VN.n181 4.5005
R11261 VN.n260 VN.n259 4.5005
R11262 VN.n262 VN.n261 4.5005
R11263 VN.n178 VN.n177 4.5005
R11264 VN.n270 VN.n269 4.5005
R11265 VN.n271 VN.n176 4.5005
R11266 VN.n273 VN.n272 4.5005
R11267 VN.n174 VN.n173 4.5005
R11268 VN.n280 VN.n279 4.5005
R11269 VN.n282 VN.n281 4.5005
R11270 VN.n170 VN.n169 4.5005
R11271 VN.n289 VN.n288 4.5005
R11272 VN.n291 VN.n290 4.5005
R11273 VN.n166 VN.n165 4.5005
R11274 VN.n298 VN.n297 4.5005
R11275 VN.n300 VN.n299 4.5005
R11276 VN.n162 VN.n161 4.5005
R11277 VN.n308 VN.n307 4.5005
R11278 VN.n309 VN.n160 4.5005
R11279 VN.n311 VN.n310 4.5005
R11280 VN.n158 VN.n157 4.5005
R11281 VN.n318 VN.n317 4.5005
R11282 VN.n376 VN.n375 4.5005
R11283 VN.n374 VN.n373 4.5005
R11284 VN.n334 VN.n332 4.5005
R11285 VN.n368 VN.n367 4.5005
R11286 VN.n366 VN.n365 4.5005
R11287 VN.n339 VN.n337 4.5005
R11288 VN.n360 VN.n359 4.5005
R11289 VN.n358 VN.n357 4.5005
R11290 VN.n344 VN.n342 4.5005
R11291 VN.n348 VN.n346 4.5005
R11292 VN.n352 VN.n351 4.5005
R11293 VN.n204 VN.n203 4.5005
R11294 VN.n206 VN.n205 4.5005
R11295 VN.n198 VN.n197 4.5005
R11296 VN.n214 VN.n213 4.5005
R11297 VN.n216 VN.n215 4.5005
R11298 VN.n218 VN.n193 4.5005
R11299 VN.n224 VN.n223 4.5005
R11300 VN.n225 VN.n192 4.5005
R11301 VN.n227 VN.n226 4.5005
R11302 VN.n229 VN.n189 4.5005
R11303 VN.n234 VN.n233 4.5005
R11304 VN.n200 VN.n199 4.5005
R11305 VN.n208 VN.n207 4.5005
R11306 VN.n211 VN.n210 4.5005
R11307 VN.n209 VN.n196 4.5005
R11308 VN.n217 VN.n195 4.5005
R11309 VN.n220 VN.n219 4.5005
R11310 VN.n222 VN.n221 4.5005
R11311 VN.n228 VN.n191 4.5005
R11312 VN.n231 VN.n230 4.5005
R11313 VN.n249 VN.n183 4.5005
R11314 VN.n255 VN.n254 4.5005
R11315 VN.n257 VN.n256 4.5005
R11316 VN.n258 VN.n179 4.5005
R11317 VN.n264 VN.n263 4.5005
R11318 VN.n266 VN.n265 4.5005
R11319 VN.n268 VN.n175 4.5005
R11320 VN.n275 VN.n274 4.5005
R11321 VN.n277 VN.n276 4.5005
R11322 VN.n278 VN.n171 4.5005
R11323 VN.n286 VN.n285 4.5005
R11324 VN.n168 VN.n167 4.5005
R11325 VN.n293 VN.n292 4.5005
R11326 VN.n295 VN.n294 4.5005
R11327 VN.n164 VN.n163 4.5005
R11328 VN.n302 VN.n301 4.5005
R11329 VN.n304 VN.n303 4.5005
R11330 VN.n306 VN.n159 4.5005
R11331 VN.n313 VN.n312 4.5005
R11332 VN.n315 VN.n314 4.5005
R11333 VN.n152 VN.n151 4.5005
R11334 VN.n372 VN.n371 4.5005
R11335 VN.n370 VN.n369 4.5005
R11336 VN.n336 VN.n335 4.5005
R11337 VN.n364 VN.n363 4.5005
R11338 VN.n362 VN.n361 4.5005
R11339 VN.n341 VN.n340 4.5005
R11340 VN.n356 VN.n355 4.5005
R11341 VN.n354 VN.n353 4.5005
R11342 VN.n347 VN.n345 4.5005
R11343 VN.n113 VN.n62 4.5005
R11344 VN.n112 VN.n111 4.5005
R11345 VN.n110 VN.n63 4.5005
R11346 VN.n109 VN.n108 4.5005
R11347 VN.n106 VN.n64 4.5005
R11348 VN.n105 VN.n104 4.5005
R11349 VN.n428 VN.n427 4.5005
R11350 VN.n429 VN.n385 4.5005
R11351 VN.n431 VN.n430 4.5005
R11352 VN.n432 VN.n384 4.5005
R11353 VN.n434 VN.n433 4.5005
R11354 VN.n435 VN.n383 4.5005
R11355 VN.n461 VN.n460 4.5005
R11356 VN.n134 VN.n131 4.5005
R11357 VN.n465 VN.n130 4.5005
R11358 VN.n466 VN.n129 4.5005
R11359 VN.n467 VN.n128 4.5005
R11360 VN.n470 VN.n125 4.5005
R11361 VN.n471 VN.n124 4.5005
R11362 VN.n472 VN.n123 4.5005
R11363 VN.n122 VN.n119 4.5005
R11364 VN.n476 VN.n118 4.5005
R11365 VN.n477 VN.n117 4.5005
R11366 VN.n479 VN.n116 4.5005
R11367 VN.n439 VN.n438 4.5005
R11368 VN.n382 VN.n149 4.5005
R11369 VN.n443 VN.n148 4.5005
R11370 VN.n444 VN.n147 4.5005
R11371 VN.n445 VN.n146 4.5005
R11372 VN.n145 VN.n142 4.5005
R11373 VN.n449 VN.n141 4.5005
R11374 VN.n450 VN.n140 4.5005
R11375 VN.n452 VN.n139 4.5005
R11376 VN.n138 VN.n136 4.5005
R11377 VN.n456 VN.n135 4.5005
R11378 VN.n459 VN.n458 4.5005
R11379 VN.n405 VN.n403 4.5005
R11380 VN.n409 VN.n402 4.5005
R11381 VN.n410 VN.n401 4.5005
R11382 VN.n411 VN.n400 4.5005
R11383 VN.n414 VN.n397 4.5005
R11384 VN.n415 VN.n396 4.5005
R11385 VN.n416 VN.n395 4.5005
R11386 VN.n419 VN.n392 4.5005
R11387 VN.n420 VN.n391 4.5005
R11388 VN.n421 VN.n388 4.5005
R11389 VN.n425 VN.n424 4.5005
R11390 VN.n102 VN.n101 4.5005
R11391 VN.n99 VN.n66 4.5005
R11392 VN.n93 VN.n67 4.5005
R11393 VN.n95 VN.n94 4.5005
R11394 VN.n92 VN.n69 4.5005
R11395 VN.n91 VN.n90 4.5005
R11396 VN.n71 VN.n70 4.5005
R11397 VN.n86 VN.n85 4.5005
R11398 VN.n84 VN.n83 4.5005
R11399 VN.n82 VN.n75 4.5005
R11400 VN.n77 VN.n76 4.5005
R11401 VN.n80 VN.n76 4.5005
R11402 VN.n82 VN.n81 4.5005
R11403 VN.n83 VN.n73 4.5005
R11404 VN.n87 VN.n86 4.5005
R11405 VN.n88 VN.n71 4.5005
R11406 VN.n90 VN.n89 4.5005
R11407 VN.n69 VN.n68 4.5005
R11408 VN.n96 VN.n95 4.5005
R11409 VN.n97 VN.n67 4.5005
R11410 VN.n99 VN.n98 4.5005
R11411 VN.n101 VN.n60 4.5005
R11412 VN.n480 VN.n479 4.5005
R11413 VN.n477 VN.n61 4.5005
R11414 VN.n476 VN.n475 4.5005
R11415 VN.n474 VN.n119 4.5005
R11416 VN.n473 VN.n472 4.5005
R11417 VN.n471 VN.n120 4.5005
R11418 VN.n470 VN.n469 4.5005
R11419 VN.n468 VN.n467 4.5005
R11420 VN.n466 VN.n127 4.5005
R11421 VN.n465 VN.n464 4.5005
R11422 VN.n463 VN.n131 4.5005
R11423 VN.n462 VN.n461 4.5005
R11424 VN.n458 VN.n132 4.5005
R11425 VN.n456 VN.n455 4.5005
R11426 VN.n454 VN.n136 4.5005
R11427 VN.n453 VN.n452 4.5005
R11428 VN.n450 VN.n137 4.5005
R11429 VN.n449 VN.n448 4.5005
R11430 VN.n447 VN.n142 4.5005
R11431 VN.n446 VN.n445 4.5005
R11432 VN.n444 VN.n143 4.5005
R11433 VN.n443 VN.n442 4.5005
R11434 VN.n441 VN.n149 4.5005
R11435 VN.n440 VN.n439 4.5005
R11436 VN.n424 VN.n423 4.5005
R11437 VN.n422 VN.n421 4.5005
R11438 VN.n420 VN.n390 4.5005
R11439 VN.n419 VN.n418 4.5005
R11440 VN.n417 VN.n416 4.5005
R11441 VN.n415 VN.n394 4.5005
R11442 VN.n414 VN.n413 4.5005
R11443 VN.n412 VN.n411 4.5005
R11444 VN.n410 VN.n399 4.5005
R11445 VN.n409 VN.n408 4.5005
R11446 VN.n407 VN.n403 4.5005
R11447 VN.n545 VN.n486 4.5005
R11448 VN.n544 VN.n543 4.5005
R11449 VN.n542 VN.n487 4.5005
R11450 VN.n541 VN.n540 4.5005
R11451 VN.n538 VN.n488 4.5005
R11452 VN.n537 VN.n536 4.5005
R11453 VN.n638 VN.n637 4.5005
R11454 VN.n639 VN.n584 4.5005
R11455 VN.n641 VN.n640 4.5005
R11456 VN.n642 VN.n583 4.5005
R11457 VN.n644 VN.n643 4.5005
R11458 VN.n645 VN.n582 4.5005
R11459 VN.n710 VN.n709 4.5005
R11460 VN.n708 VN.n707 4.5005
R11461 VN.n550 VN.n548 4.5005
R11462 VN.n702 VN.n701 4.5005
R11463 VN.n700 VN.n699 4.5005
R11464 VN.n555 VN.n553 4.5005
R11465 VN.n694 VN.n693 4.5005
R11466 VN.n692 VN.n691 4.5005
R11467 VN.n560 VN.n558 4.5005
R11468 VN.n564 VN.n562 4.5005
R11469 VN.n686 VN.n685 4.5005
R11470 VN.n684 VN.n683 4.5005
R11471 VN.n680 VN.n565 4.5005
R11472 VN.n677 VN.n676 4.5005
R11473 VN.n675 VN.n674 4.5005
R11474 VN.n570 VN.n569 4.5005
R11475 VN.n668 VN.n667 4.5005
R11476 VN.n666 VN.n665 4.5005
R11477 VN.n575 VN.n574 4.5005
R11478 VN.n659 VN.n658 4.5005
R11479 VN.n657 VN.n656 4.5005
R11480 VN.n655 VN.n578 4.5005
R11481 VN.n581 VN.n579 4.5005
R11482 VN.n649 VN.n648 4.5005
R11483 VN.n635 VN.n634 4.5005
R11484 VN.n592 VN.n587 4.5005
R11485 VN.n629 VN.n628 4.5005
R11486 VN.n627 VN.n626 4.5005
R11487 VN.n597 VN.n594 4.5005
R11488 VN.n621 VN.n620 4.5005
R11489 VN.n619 VN.n618 4.5005
R11490 VN.n602 VN.n599 4.5005
R11491 VN.n613 VN.n612 4.5005
R11492 VN.n611 VN.n603 4.5005
R11493 VN.n610 VN.n609 4.5005
R11494 VN.n505 VN.n504 4.5005
R11495 VN.n507 VN.n506 4.5005
R11496 VN.n499 VN.n498 4.5005
R11497 VN.n514 VN.n513 4.5005
R11498 VN.n516 VN.n515 4.5005
R11499 VN.n495 VN.n494 4.5005
R11500 VN.n524 VN.n523 4.5005
R11501 VN.n525 VN.n493 4.5005
R11502 VN.n527 VN.n526 4.5005
R11503 VN.n491 VN.n490 4.5005
R11504 VN.n534 VN.n533 4.5005
R11505 VN.n501 VN.n500 4.5005
R11506 VN.n509 VN.n508 4.5005
R11507 VN.n511 VN.n510 4.5005
R11508 VN.n497 VN.n496 4.5005
R11509 VN.n518 VN.n517 4.5005
R11510 VN.n520 VN.n519 4.5005
R11511 VN.n522 VN.n492 4.5005
R11512 VN.n529 VN.n528 4.5005
R11513 VN.n531 VN.n530 4.5005
R11514 VN.n485 VN.n484 4.5005
R11515 VN.n706 VN.n705 4.5005
R11516 VN.n704 VN.n703 4.5005
R11517 VN.n552 VN.n551 4.5005
R11518 VN.n698 VN.n697 4.5005
R11519 VN.n696 VN.n695 4.5005
R11520 VN.n557 VN.n556 4.5005
R11521 VN.n690 VN.n689 4.5005
R11522 VN.n688 VN.n687 4.5005
R11523 VN.n563 VN.n561 4.5005
R11524 VN.n679 VN.n567 4.5005
R11525 VN.n571 VN.n568 4.5005
R11526 VN.n673 VN.n672 4.5005
R11527 VN.n671 VN.n670 4.5005
R11528 VN.n573 VN.n572 4.5005
R11529 VN.n664 VN.n663 4.5005
R11530 VN.n662 VN.n661 4.5005
R11531 VN.n577 VN.n576 4.5005
R11532 VN.n654 VN.n653 4.5005
R11533 VN.n652 VN.n651 4.5005
R11534 VN.n633 VN.n632 4.5005
R11535 VN.n631 VN.n630 4.5005
R11536 VN.n593 VN.n591 4.5005
R11537 VN.n625 VN.n624 4.5005
R11538 VN.n623 VN.n622 4.5005
R11539 VN.n598 VN.n596 4.5005
R11540 VN.n617 VN.n616 4.5005
R11541 VN.n615 VN.n614 4.5005
R11542 VN.n605 VN.n601 4.5005
R11543 VN.n608 VN.n607 4.5005
R11544 VN.n843 VN.n842 4.5005
R11545 VN.n840 VN.n715 4.5005
R11546 VN.n773 VN.n771 4.5005
R11547 VN.n836 VN.n774 4.5005
R11548 VN.n834 VN.n775 4.5005
R11549 VN.n833 VN.n776 4.5005
R11550 VN.n780 VN.n777 4.5005
R11551 VN.n829 VN.n781 4.5005
R11552 VN.n828 VN.n782 4.5005
R11553 VN.n827 VN.n783 4.5005
R11554 VN.n787 VN.n784 4.5005
R11555 VN.n823 VN.n822 4.5005
R11556 VN.n57 VN.n56 4.5005
R11557 VN.n54 VN.n3 4.5005
R11558 VN.n24 VN.n22 4.5005
R11559 VN.n50 VN.n25 4.5005
R11560 VN.n48 VN.n26 4.5005
R11561 VN.n47 VN.n27 4.5005
R11562 VN.n31 VN.n28 4.5005
R11563 VN.n43 VN.n32 4.5005
R11564 VN.n42 VN.n33 4.5005
R11565 VN.n41 VN.n34 4.5005
R11566 VN.n37 VN.n35 4.5005
R11567 VN.n733 VN.n729 4.5005
R11568 VN.n735 VN.n734 4.5005
R11569 VN.n736 VN.n726 4.5005
R11570 VN.n740 VN.n739 4.5005
R11571 VN.n741 VN.n725 4.5005
R11572 VN.n744 VN.n742 4.5005
R11573 VN.n723 VN.n722 4.5005
R11574 VN.n750 VN.n749 4.5005
R11575 VN.n751 VN.n721 4.5005
R11576 VN.n753 VN.n752 4.5005
R11577 VN.n755 VN.n714 4.5005
R11578 VN.n767 VN.n716 4.5005
R11579 VN.n766 VN.n765 4.5005
R11580 VN.n764 VN.n717 4.5005
R11581 VN.n763 VN.n762 4.5005
R11582 VN.n760 VN.n718 4.5005
R11583 VN.n759 VN.n758 4.5005
R11584 VN.n18 VN.n4 4.5005
R11585 VN.n17 VN.n16 4.5005
R11586 VN.n15 VN.n5 4.5005
R11587 VN.n14 VN.n13 4.5005
R11588 VN.n11 VN.n6 4.5005
R11589 VN.n10 VN.n9 4.5005
R11590 VN.n756 VN.n755 4.5005
R11591 VN.n753 VN.n720 4.5005
R11592 VN.n747 VN.n721 4.5005
R11593 VN.n749 VN.n748 4.5005
R11594 VN.n746 VN.n723 4.5005
R11595 VN.n745 VN.n744 4.5005
R11596 VN.n725 VN.n724 4.5005
R11597 VN.n739 VN.n738 4.5005
R11598 VN.n737 VN.n736 4.5005
R11599 VN.n735 VN.n728 4.5005
R11600 VN.n731 VN.n729 4.5005
R11601 VN.n824 VN.n823 4.5005
R11602 VN.n825 VN.n784 4.5005
R11603 VN.n827 VN.n826 4.5005
R11604 VN.n828 VN.n778 4.5005
R11605 VN.n830 VN.n829 4.5005
R11606 VN.n831 VN.n777 4.5005
R11607 VN.n833 VN.n832 4.5005
R11608 VN.n834 VN.n772 4.5005
R11609 VN.n837 VN.n836 4.5005
R11610 VN.n838 VN.n771 4.5005
R11611 VN.n840 VN.n839 4.5005
R11612 VN.n842 VN.n770 4.5005
R11613 VN.n39 VN.n35 4.5005
R11614 VN.n41 VN.n40 4.5005
R11615 VN.n42 VN.n29 4.5005
R11616 VN.n44 VN.n43 4.5005
R11617 VN.n45 VN.n28 4.5005
R11618 VN.n47 VN.n46 4.5005
R11619 VN.n48 VN.n23 4.5005
R11620 VN.n51 VN.n50 4.5005
R11621 VN.n52 VN.n22 4.5005
R11622 VN.n54 VN.n53 4.5005
R11623 VN.n56 VN.n21 4.5005
R11624 VN.n849 VN.n1 4.5005
R11625 VN.n804 VN.n803 4.5005
R11626 VN.n806 VN.n802 4.5005
R11627 VN.n807 VN.n801 4.5005
R11628 VN.n808 VN.n800 4.5005
R11629 VN.n811 VN.n797 4.5005
R11630 VN.n812 VN.n796 4.5005
R11631 VN.n813 VN.n795 4.5005
R11632 VN.n794 VN.n791 4.5005
R11633 VN.n817 VN.n790 4.5005
R11634 VN.n818 VN.n789 4.5005
R11635 VN.n820 VN.n785 4.5005
R11636 VN.n821 VN.n820 4.5005
R11637 VN.n818 VN.n788 4.5005
R11638 VN.n817 VN.n816 4.5005
R11639 VN.n815 VN.n791 4.5005
R11640 VN.n814 VN.n813 4.5005
R11641 VN.n812 VN.n792 4.5005
R11642 VN.n811 VN.n810 4.5005
R11643 VN.n809 VN.n808 4.5005
R11644 VN.n807 VN.n799 4.5005
R11645 VN.n806 VN.n805 4.5005
R11646 VN.n804 VN.n2 4.5005
R11647 VN.n849 VN.n848 4.5005
R11648 VN.n281 VN.n169 3.0245
R11649 VN.n460 VN.n459 3.0245
R11650 VN.n462 VN.n132 3.0245
R11651 VN.n684 VN.n565 3.0245
R11652 VN.n822 VN.n821 3.0245
R11653 VN.n824 VN.n785 3.0245
R11654 VN.n284 VN.n283 2.96825
R11655 VN.n682 VN.n681 2.96825
R11656 VN.n201 VN.n199 2.41967
R11657 VN.n502 VN.n500 2.41967
R11658 VN.n437 VN.n436 2.22849
R11659 VN.n103 VN.n65 2.22849
R11660 VN.n8 VN.n7 2.22849
R11661 VN.n757 VN.n719 2.22849
R11662 VN.n319 VN.n156 2.22782
R11663 VN.n235 VN.n188 2.22782
R11664 VN.n647 VN.n646 2.22782
R11665 VN.n535 VN.n489 2.22782
R11666 VN.n481 VN.n480 2.102
R11667 VN.n423 VN.n380 2.102
R11668 VN.n844 VN.n843 2.102
R11669 VN.n847 VN.n57 2.102
R11670 VN.n482 VN.n59 2.07182
R11671 VN.n379 VN.n378 2.07182
R11672 VN.n248 VN.n59 2.06825
R11673 VN.n378 VN.n377 2.06825
R11674 VN.n712 VN.n711 2.06825
R11675 VN.n589 VN.n588 2.06825
R11676 VN.n713 VN.n712 1.5005
R11677 VN.n482 VN.n481 1.5005
R11678 VN.n588 VN.n58 1.5005
R11679 VN.n380 VN.n379 1.5005
R11680 VN.n847 VN.n846 1.5005
R11681 VN.n845 VN.n844 1.5005
R11682 VN.n713 VN.n482 1.47516
R11683 VN.n379 VN.n58 1.47516
R11684 VN.n481 VN.n60 0.83975
R11685 VN.n440 VN.n380 0.83975
R11686 VN.n844 VN.n714 0.83975
R11687 VN.n848 VN.n847 0.83975
R11688 VN.n232 VN.n59 0.81725
R11689 VN.n378 VN.n150 0.81725
R11690 VN.n712 VN.n483 0.81725
R11691 VN.n588 VN.n580 0.81725
R11692 VN.n103 VN.n102 0.75626
R11693 VN.n438 VN.n437 0.75626
R11694 VN.n757 VN.n756 0.75626
R11695 VN.n8 VN.n1 0.75626
R11696 VN.n235 VN.n234 0.756242
R11697 VN.n319 VN.n318 0.756242
R11698 VN.n535 VN.n534 0.756242
R11699 VN.n648 VN.n647 0.756242
R11700 VN.n251 VN.n247 0.698
R11701 VN.n375 VN.n331 0.698
R11702 VN.n116 VN.n115 0.698
R11703 VN.n426 VN.n425 0.698
R11704 VN.n709 VN.n547 0.698
R11705 VN.n636 VN.n635 0.698
R11706 VN.n770 VN.n769 0.698
R11707 VN.n21 VN.n20 0.698
R11708 VN.n845 VN.n713 0.571818
R11709 VN.n846 VN.n58 0.571818
R11710 VN.n215 VN.n193 0.375125
R11711 VN.n270 VN.n177 0.375125
R11712 VN.n299 VN.n161 0.375125
R11713 VN.n359 VN.n337 0.375125
R11714 VN.n91 VN.n70 0.375125
R11715 VN.n125 VN.n124 0.375125
R11716 VN.n145 VN.n141 0.375125
R11717 VN.n397 VN.n396 0.375125
R11718 VN.n89 VN.n88 0.375125
R11719 VN.n469 VN.n120 0.375125
R11720 VN.n448 VN.n447 0.375125
R11721 VN.n413 VN.n394 0.375125
R11722 VN.n515 VN.n494 0.375125
R11723 VN.n693 VN.n553 0.375125
R11724 VN.n666 VN.n574 0.375125
R11725 VN.n620 VN.n619 0.375125
R11726 VN.n742 VN.n741 0.375125
R11727 VN.n780 VN.n776 0.375125
R11728 VN.n810 VN.n792 0.375125
R11729 VN.n31 VN.n27 0.375125
R11730 VN.n745 VN.n724 0.375125
R11731 VN.n832 VN.n831 0.375125
R11732 VN.n797 VN.n796 0.375125
R11733 VN.n46 VN.n45 0.375125
R11734 VN.n205 VN.n197 0.36275
R11735 VN.n260 VN.n181 0.36275
R11736 VN.n290 VN.n165 0.36275
R11737 VN.n367 VN.n332 0.36275
R11738 VN.n84 VN.n75 0.36275
R11739 VN.n122 VN.n118 0.36275
R11740 VN.n139 VN.n138 0.36275
R11741 VN.n392 VN.n391 0.36275
R11742 VN.n81 VN.n73 0.36275
R11743 VN.n475 VN.n474 0.36275
R11744 VN.n454 VN.n453 0.36275
R11745 VN.n418 VN.n390 0.36275
R11746 VN.n506 VN.n498 0.36275
R11747 VN.n701 VN.n548 0.36275
R11748 VN.n675 VN.n569 0.36275
R11749 VN.n628 VN.n627 0.36275
R11750 VN.n734 VN.n726 0.36275
R11751 VN.n774 VN.n773 0.36275
R11752 VN.n816 VN.n815 0.36275
R11753 VN.n25 VN.n24 0.36275
R11754 VN.n737 VN.n728 0.36275
R11755 VN.n838 VN.n837 0.36275
R11756 VN.n794 VN.n790 0.36275
R11757 VN.n52 VN.n51 0.36275
R11758 VN.n236 VN.n187 0.3605
R11759 VN.n243 VN.n242 0.3605
R11760 VN.n320 VN.n155 0.3605
R11761 VN.n327 VN.n326 0.3605
R11762 VN.n208 VN.n199 0.3605
R11763 VN.n209 VN.n195 0.3605
R11764 VN.n221 VN.n191 0.3605
R11765 VN.n256 VN.n255 0.3605
R11766 VN.n265 VN.n264 0.3605
R11767 VN.n276 VN.n275 0.3605
R11768 VN.n293 VN.n167 0.3605
R11769 VN.n302 VN.n163 0.3605
R11770 VN.n313 VN.n159 0.3605
R11771 VN.n371 VN.n370 0.3605
R11772 VN.n363 VN.n362 0.3605
R11773 VN.n355 VN.n354 0.3605
R11774 VN.n104 VN.n64 0.3605
R11775 VN.n111 VN.n110 0.3605
R11776 VN.n433 VN.n383 0.3605
R11777 VN.n431 VN.n385 0.3605
R11778 VN.n536 VN.n488 0.3605
R11779 VN.n543 VN.n542 0.3605
R11780 VN.n643 VN.n582 0.3605
R11781 VN.n641 VN.n584 0.3605
R11782 VN.n509 VN.n500 0.3605
R11783 VN.n518 VN.n496 0.3605
R11784 VN.n529 VN.n492 0.3605
R11785 VN.n705 VN.n704 0.3605
R11786 VN.n697 VN.n696 0.3605
R11787 VN.n689 VN.n688 0.3605
R11788 VN.n672 VN.n571 0.3605
R11789 VN.n663 VN.n572 0.3605
R11790 VN.n653 VN.n576 0.3605
R11791 VN.n631 VN.n591 0.3605
R11792 VN.n623 VN.n596 0.3605
R11793 VN.n615 VN.n601 0.3605
R11794 VN.n758 VN.n718 0.3605
R11795 VN.n765 VN.n764 0.3605
R11796 VN.n9 VN.n6 0.3605
R11797 VN.n16 VN.n15 0.3605
R11798 VN.n226 VN.n225 0.287375
R11799 VN.n272 VN.n173 0.287375
R11800 VN.n310 VN.n309 0.287375
R11801 VN.n348 VN.n342 0.287375
R11802 VN.n94 VN.n93 0.287375
R11803 VN.n130 VN.n129 0.287375
R11804 VN.n148 VN.n147 0.287375
R11805 VN.n402 VN.n401 0.287375
R11806 VN.n97 VN.n96 0.287375
R11807 VN.n464 VN.n127 0.287375
R11808 VN.n442 VN.n143 0.287375
R11809 VN.n408 VN.n399 0.287375
R11810 VN.n526 VN.n525 0.287375
R11811 VN.n564 VN.n558 0.287375
R11812 VN.n657 VN.n578 0.287375
R11813 VN.n612 VN.n611 0.287375
R11814 VN.n751 VN.n750 0.287375
R11815 VN.n783 VN.n782 0.287375
R11816 VN.n805 VN.n799 0.287375
R11817 VN.n34 VN.n33 0.287375
R11818 VN.n748 VN.n747 0.287375
R11819 VN.n826 VN.n778 0.287375
R11820 VN.n802 VN.n801 0.287375
R11821 VN.n40 VN.n29 0.287375
R11822 VN.n236 VN.n235 0.208888
R11823 VN.n320 VN.n319 0.208888
R11824 VN.n536 VN.n535 0.208888
R11825 VN.n647 VN.n582 0.208888
R11826 VN.n104 VN.n103 0.20887
R11827 VN.n437 VN.n383 0.20887
R11828 VN.n758 VN.n757 0.20887
R11829 VN.n9 VN.n8 0.20887
R11830 VN.n205 VN.n204 0.14
R11831 VN.n214 VN.n197 0.14
R11832 VN.n215 VN.n214 0.14
R11833 VN.n224 VN.n193 0.14
R11834 VN.n225 VN.n224 0.14
R11835 VN.n226 VN.n189 0.14
R11836 VN.n234 VN.n189 0.14
R11837 VN.n241 VN.n187 0.14
R11838 VN.n242 VN.n241 0.14
R11839 VN.n243 VN.n185 0.14
R11840 VN.n247 VN.n185 0.14
R11841 VN.n252 VN.n251 0.14
R11842 VN.n252 VN.n181 0.14
R11843 VN.n261 VN.n260 0.14
R11844 VN.n261 VN.n177 0.14
R11845 VN.n271 VN.n270 0.14
R11846 VN.n272 VN.n271 0.14
R11847 VN.n280 VN.n173 0.14
R11848 VN.n281 VN.n280 0.14
R11849 VN.n289 VN.n169 0.14
R11850 VN.n290 VN.n289 0.14
R11851 VN.n298 VN.n165 0.14
R11852 VN.n299 VN.n298 0.14
R11853 VN.n308 VN.n161 0.14
R11854 VN.n309 VN.n308 0.14
R11855 VN.n310 VN.n157 0.14
R11856 VN.n318 VN.n157 0.14
R11857 VN.n325 VN.n155 0.14
R11858 VN.n326 VN.n325 0.14
R11859 VN.n327 VN.n153 0.14
R11860 VN.n331 VN.n153 0.14
R11861 VN.n375 VN.n374 0.14
R11862 VN.n374 VN.n332 0.14
R11863 VN.n367 VN.n366 0.14
R11864 VN.n366 VN.n337 0.14
R11865 VN.n359 VN.n358 0.14
R11866 VN.n358 VN.n342 0.14
R11867 VN.n351 VN.n348 0.14
R11868 VN.n210 VN.n208 0.14
R11869 VN.n210 VN.n209 0.14
R11870 VN.n220 VN.n195 0.14
R11871 VN.n221 VN.n220 0.14
R11872 VN.n231 VN.n191 0.14
R11873 VN.n232 VN.n231 0.14
R11874 VN.n248 VN.n183 0.14
R11875 VN.n255 VN.n183 0.14
R11876 VN.n256 VN.n179 0.14
R11877 VN.n264 VN.n179 0.14
R11878 VN.n265 VN.n175 0.14
R11879 VN.n275 VN.n175 0.14
R11880 VN.n276 VN.n171 0.14
R11881 VN.n283 VN.n171 0.14
R11882 VN.n285 VN.n284 0.14
R11883 VN.n285 VN.n167 0.14
R11884 VN.n294 VN.n293 0.14
R11885 VN.n294 VN.n163 0.14
R11886 VN.n303 VN.n302 0.14
R11887 VN.n303 VN.n159 0.14
R11888 VN.n314 VN.n313 0.14
R11889 VN.n314 VN.n150 0.14
R11890 VN.n377 VN.n151 0.14
R11891 VN.n371 VN.n151 0.14
R11892 VN.n370 VN.n335 0.14
R11893 VN.n363 VN.n335 0.14
R11894 VN.n362 VN.n340 0.14
R11895 VN.n355 VN.n340 0.14
R11896 VN.n354 VN.n345 0.14
R11897 VN.n77 VN.n75 0.14
R11898 VN.n85 VN.n84 0.14
R11899 VN.n85 VN.n70 0.14
R11900 VN.n92 VN.n91 0.14
R11901 VN.n94 VN.n92 0.14
R11902 VN.n93 VN.n66 0.14
R11903 VN.n102 VN.n66 0.14
R11904 VN.n109 VN.n64 0.14
R11905 VN.n110 VN.n109 0.14
R11906 VN.n111 VN.n62 0.14
R11907 VN.n115 VN.n62 0.14
R11908 VN.n117 VN.n116 0.14
R11909 VN.n118 VN.n117 0.14
R11910 VN.n123 VN.n122 0.14
R11911 VN.n124 VN.n123 0.14
R11912 VN.n128 VN.n125 0.14
R11913 VN.n129 VN.n128 0.14
R11914 VN.n134 VN.n130 0.14
R11915 VN.n460 VN.n134 0.14
R11916 VN.n459 VN.n135 0.14
R11917 VN.n138 VN.n135 0.14
R11918 VN.n140 VN.n139 0.14
R11919 VN.n141 VN.n140 0.14
R11920 VN.n146 VN.n145 0.14
R11921 VN.n147 VN.n146 0.14
R11922 VN.n382 VN.n148 0.14
R11923 VN.n438 VN.n382 0.14
R11924 VN.n433 VN.n432 0.14
R11925 VN.n432 VN.n431 0.14
R11926 VN.n427 VN.n385 0.14
R11927 VN.n427 VN.n426 0.14
R11928 VN.n425 VN.n388 0.14
R11929 VN.n391 VN.n388 0.14
R11930 VN.n395 VN.n392 0.14
R11931 VN.n396 VN.n395 0.14
R11932 VN.n400 VN.n397 0.14
R11933 VN.n401 VN.n400 0.14
R11934 VN.n405 VN.n402 0.14
R11935 VN.n81 VN.n80 0.14
R11936 VN.n87 VN.n73 0.14
R11937 VN.n88 VN.n87 0.14
R11938 VN.n89 VN.n68 0.14
R11939 VN.n96 VN.n68 0.14
R11940 VN.n98 VN.n97 0.14
R11941 VN.n98 VN.n60 0.14
R11942 VN.n480 VN.n61 0.14
R11943 VN.n475 VN.n61 0.14
R11944 VN.n474 VN.n473 0.14
R11945 VN.n473 VN.n120 0.14
R11946 VN.n469 VN.n468 0.14
R11947 VN.n468 VN.n127 0.14
R11948 VN.n464 VN.n463 0.14
R11949 VN.n463 VN.n462 0.14
R11950 VN.n455 VN.n132 0.14
R11951 VN.n455 VN.n454 0.14
R11952 VN.n453 VN.n137 0.14
R11953 VN.n448 VN.n137 0.14
R11954 VN.n447 VN.n446 0.14
R11955 VN.n446 VN.n143 0.14
R11956 VN.n442 VN.n441 0.14
R11957 VN.n441 VN.n440 0.14
R11958 VN.n423 VN.n422 0.14
R11959 VN.n422 VN.n390 0.14
R11960 VN.n418 VN.n417 0.14
R11961 VN.n417 VN.n394 0.14
R11962 VN.n413 VN.n412 0.14
R11963 VN.n412 VN.n399 0.14
R11964 VN.n408 VN.n407 0.14
R11965 VN.n506 VN.n505 0.14
R11966 VN.n514 VN.n498 0.14
R11967 VN.n515 VN.n514 0.14
R11968 VN.n524 VN.n494 0.14
R11969 VN.n525 VN.n524 0.14
R11970 VN.n526 VN.n490 0.14
R11971 VN.n534 VN.n490 0.14
R11972 VN.n541 VN.n488 0.14
R11973 VN.n542 VN.n541 0.14
R11974 VN.n543 VN.n486 0.14
R11975 VN.n547 VN.n486 0.14
R11976 VN.n709 VN.n708 0.14
R11977 VN.n708 VN.n548 0.14
R11978 VN.n701 VN.n700 0.14
R11979 VN.n700 VN.n553 0.14
R11980 VN.n693 VN.n692 0.14
R11981 VN.n692 VN.n558 0.14
R11982 VN.n685 VN.n564 0.14
R11983 VN.n685 VN.n684 0.14
R11984 VN.n676 VN.n565 0.14
R11985 VN.n676 VN.n675 0.14
R11986 VN.n667 VN.n569 0.14
R11987 VN.n667 VN.n666 0.14
R11988 VN.n658 VN.n574 0.14
R11989 VN.n658 VN.n657 0.14
R11990 VN.n581 VN.n578 0.14
R11991 VN.n648 VN.n581 0.14
R11992 VN.n643 VN.n642 0.14
R11993 VN.n642 VN.n641 0.14
R11994 VN.n637 VN.n584 0.14
R11995 VN.n637 VN.n636 0.14
R11996 VN.n635 VN.n587 0.14
R11997 VN.n628 VN.n587 0.14
R11998 VN.n627 VN.n594 0.14
R11999 VN.n620 VN.n594 0.14
R12000 VN.n619 VN.n599 0.14
R12001 VN.n612 VN.n599 0.14
R12002 VN.n611 VN.n610 0.14
R12003 VN.n510 VN.n509 0.14
R12004 VN.n510 VN.n496 0.14
R12005 VN.n519 VN.n518 0.14
R12006 VN.n519 VN.n492 0.14
R12007 VN.n530 VN.n529 0.14
R12008 VN.n530 VN.n483 0.14
R12009 VN.n711 VN.n484 0.14
R12010 VN.n705 VN.n484 0.14
R12011 VN.n704 VN.n551 0.14
R12012 VN.n697 VN.n551 0.14
R12013 VN.n696 VN.n556 0.14
R12014 VN.n689 VN.n556 0.14
R12015 VN.n688 VN.n561 0.14
R12016 VN.n682 VN.n561 0.14
R12017 VN.n681 VN.n567 0.14
R12018 VN.n571 VN.n567 0.14
R12019 VN.n672 VN.n671 0.14
R12020 VN.n671 VN.n572 0.14
R12021 VN.n663 VN.n662 0.14
R12022 VN.n662 VN.n576 0.14
R12023 VN.n653 VN.n652 0.14
R12024 VN.n652 VN.n580 0.14
R12025 VN.n632 VN.n589 0.14
R12026 VN.n632 VN.n631 0.14
R12027 VN.n624 VN.n591 0.14
R12028 VN.n624 VN.n623 0.14
R12029 VN.n616 VN.n596 0.14
R12030 VN.n616 VN.n615 0.14
R12031 VN.n607 VN.n601 0.14
R12032 VN.n734 VN.n733 0.14
R12033 VN.n740 VN.n726 0.14
R12034 VN.n741 VN.n740 0.14
R12035 VN.n742 VN.n722 0.14
R12036 VN.n750 VN.n722 0.14
R12037 VN.n752 VN.n751 0.14
R12038 VN.n752 VN.n714 0.14
R12039 VN.n843 VN.n715 0.14
R12040 VN.n773 VN.n715 0.14
R12041 VN.n775 VN.n774 0.14
R12042 VN.n776 VN.n775 0.14
R12043 VN.n781 VN.n780 0.14
R12044 VN.n782 VN.n781 0.14
R12045 VN.n787 VN.n783 0.14
R12046 VN.n822 VN.n787 0.14
R12047 VN.n821 VN.n788 0.14
R12048 VN.n816 VN.n788 0.14
R12049 VN.n815 VN.n814 0.14
R12050 VN.n814 VN.n792 0.14
R12051 VN.n810 VN.n809 0.14
R12052 VN.n809 VN.n799 0.14
R12053 VN.n805 VN.n2 0.14
R12054 VN.n848 VN.n2 0.14
R12055 VN.n57 VN.n3 0.14
R12056 VN.n24 VN.n3 0.14
R12057 VN.n26 VN.n25 0.14
R12058 VN.n27 VN.n26 0.14
R12059 VN.n32 VN.n31 0.14
R12060 VN.n33 VN.n32 0.14
R12061 VN.n37 VN.n34 0.14
R12062 VN.n731 VN.n728 0.14
R12063 VN.n738 VN.n737 0.14
R12064 VN.n738 VN.n724 0.14
R12065 VN.n746 VN.n745 0.14
R12066 VN.n748 VN.n746 0.14
R12067 VN.n747 VN.n720 0.14
R12068 VN.n756 VN.n720 0.14
R12069 VN.n763 VN.n718 0.14
R12070 VN.n764 VN.n763 0.14
R12071 VN.n765 VN.n716 0.14
R12072 VN.n769 VN.n716 0.14
R12073 VN.n839 VN.n770 0.14
R12074 VN.n839 VN.n838 0.14
R12075 VN.n837 VN.n772 0.14
R12076 VN.n832 VN.n772 0.14
R12077 VN.n831 VN.n830 0.14
R12078 VN.n830 VN.n778 0.14
R12079 VN.n826 VN.n825 0.14
R12080 VN.n825 VN.n824 0.14
R12081 VN.n789 VN.n785 0.14
R12082 VN.n790 VN.n789 0.14
R12083 VN.n795 VN.n794 0.14
R12084 VN.n796 VN.n795 0.14
R12085 VN.n800 VN.n797 0.14
R12086 VN.n801 VN.n800 0.14
R12087 VN.n803 VN.n802 0.14
R12088 VN.n803 VN.n1 0.14
R12089 VN.n14 VN.n6 0.14
R12090 VN.n15 VN.n14 0.14
R12091 VN.n16 VN.n4 0.14
R12092 VN.n20 VN.n4 0.14
R12093 VN.n53 VN.n21 0.14
R12094 VN.n53 VN.n52 0.14
R12095 VN.n51 VN.n23 0.14
R12096 VN.n46 VN.n23 0.14
R12097 VN.n45 VN.n44 0.14
R12098 VN.n44 VN.n29 0.14
R12099 VN.n40 VN.n39 0.14
R12100 VN.n435 VN.n434 0.109179
R12101 VN.n430 VN.n429 0.109179
R12102 VN.n106 VN.n105 0.109179
R12103 VN.n112 VN.n63 0.109179
R12104 VN.n11 VN.n10 0.109179
R12105 VN.n17 VN.n5 0.109179
R12106 VN.n760 VN.n759 0.109179
R12107 VN.n766 VN.n717 0.109179
R12108 VN.n47 VN.n28 0.107155
R12109 VN.n833 VN.n777 0.107155
R12110 VN.n415 VN.n414 0.107155
R12111 VN.n449 VN.n142 0.107155
R12112 VN.n471 VN.n470 0.107155
R12113 VN.n90 VN.n71 0.107155
R12114 VN.n744 VN.n725 0.107155
R12115 VN.n812 VN.n811 0.107155
R12116 VN.n50 VN.n22 0.103632
R12117 VN.n836 VN.n771 0.103632
R12118 VN.n420 VN.n419 0.103632
R12119 VN.n452 VN.n136 0.103632
R12120 VN.n476 VN.n119 0.103632
R12121 VN.n83 VN.n82 0.103632
R12122 VN.n736 VN.n735 0.103632
R12123 VN.n817 VN.n791 0.103632
R12124 VN.n322 VN.n321 0.102991
R12125 VN.n328 VN.n154 0.102991
R12126 VN.n238 VN.n237 0.102991
R12127 VN.n244 VN.n186 0.102991
R12128 VN.n645 VN.n644 0.102991
R12129 VN.n640 VN.n639 0.102991
R12130 VN.n538 VN.n537 0.102991
R12131 VN.n544 VN.n487 0.102991
R12132 VN.n369 VN.n334 0.0933826
R12133 VN.n292 VN.n291 0.0933826
R12134 VN.n257 VN.n182 0.0933826
R12135 VN.n207 VN.n206 0.0933826
R12136 VN.n629 VN.n593 0.0933826
R12137 VN.n674 VN.n673 0.0933826
R12138 VN.n703 VN.n550 0.0933826
R12139 VN.n508 VN.n507 0.0933826
R12140 VN.n361 VN.n339 0.092742
R12141 VN.n301 VN.n300 0.092742
R12142 VN.n266 VN.n178 0.092742
R12143 VN.n217 VN.n216 0.092742
R12144 VN.n621 VN.n598 0.092742
R12145 VN.n665 VN.n664 0.092742
R12146 VN.n695 VN.n555 0.092742
R12147 VN.n517 VN.n516 0.092742
R12148 VN.n42 VN.n41 0.0821726
R12149 VN.n828 VN.n827 0.0821726
R12150 VN.n346 VN.n344 0.0821726
R12151 VN.n311 VN.n160 0.0821726
R12152 VN.n273 VN.n174 0.0821726
R12153 VN.n227 VN.n192 0.0821726
R12154 VN.n410 VN.n409 0.0821726
R12155 VN.n444 VN.n443 0.0821726
R12156 VN.n466 VN.n465 0.0821726
R12157 VN.n95 VN.n67 0.0821726
R12158 VN.n613 VN.n603 0.0821726
R12159 VN.n656 VN.n655 0.0821726
R12160 VN.n562 VN.n560 0.0821726
R12161 VN.n527 VN.n493 0.0821726
R12162 VN.n749 VN.n721 0.0821726
R12163 VN.n807 VN.n806 0.0821726
R12164 VN.n434 VN.n384 0.0426132
R12165 VN.n429 VN.n428 0.0426132
R12166 VN.n108 VN.n106 0.0426132
R12167 VN.n113 VN.n112 0.0426132
R12168 VN.n13 VN.n11 0.0426132
R12169 VN.n18 VN.n17 0.0426132
R12170 VN.n762 VN.n760 0.0426132
R12171 VN.n767 VN.n766 0.0426132
R12172 VN.n436 VN.n435 0.0412547
R12173 VN.n430 VN.n386 0.0412547
R12174 VN.n105 VN.n65 0.0412547
R12175 VN.n107 VN.n63 0.0412547
R12176 VN.n10 VN.n7 0.0412547
R12177 VN.n12 VN.n5 0.0412547
R12178 VN.n759 VN.n719 0.0412547
R12179 VN.n761 VN.n717 0.0412547
R12180 VN.n54 VN.n22 0.0402153
R12181 VN.n48 VN.n47 0.0402153
R12182 VN.n43 VN.n42 0.0402153
R12183 VN.n41 VN.n35 0.0402153
R12184 VN.n840 VN.n771 0.0402153
R12185 VN.n834 VN.n833 0.0402153
R12186 VN.n829 VN.n828 0.0402153
R12187 VN.n827 VN.n784 0.0402153
R12188 VN.n324 VN.n322 0.0402153
R12189 VN.n329 VN.n328 0.0402153
R12190 VN.n240 VN.n238 0.0402153
R12191 VN.n245 VN.n244 0.0402153
R12192 VN.n421 VN.n420 0.0402153
R12193 VN.n416 VN.n415 0.0402153
R12194 VN.n411 VN.n410 0.0402153
R12195 VN.n409 VN.n403 0.0402153
R12196 VN.n456 VN.n136 0.0402153
R12197 VN.n450 VN.n449 0.0402153
R12198 VN.n445 VN.n444 0.0402153
R12199 VN.n443 VN.n149 0.0402153
R12200 VN.n477 VN.n476 0.0402153
R12201 VN.n472 VN.n471 0.0402153
R12202 VN.n467 VN.n466 0.0402153
R12203 VN.n465 VN.n131 0.0402153
R12204 VN.n82 VN.n76 0.0402153
R12205 VN.n86 VN.n71 0.0402153
R12206 VN.n95 VN.n69 0.0402153
R12207 VN.n99 VN.n67 0.0402153
R12208 VN.n644 VN.n583 0.0402153
R12209 VN.n639 VN.n638 0.0402153
R12210 VN.n540 VN.n538 0.0402153
R12211 VN.n545 VN.n544 0.0402153
R12212 VN.n735 VN.n729 0.0402153
R12213 VN.n739 VN.n725 0.0402153
R12214 VN.n749 VN.n723 0.0402153
R12215 VN.n753 VN.n721 0.0402153
R12216 VN.n818 VN.n817 0.0402153
R12217 VN.n813 VN.n812 0.0402153
R12218 VN.n808 VN.n807 0.0402153
R12219 VN.n806 VN.n804 0.0402153
R12220 VN.n321 VN.n156 0.0389342
R12221 VN.n323 VN.n154 0.0389342
R12222 VN.n237 VN.n188 0.0389342
R12223 VN.n239 VN.n186 0.0389342
R12224 VN.n646 VN.n645 0.0389342
R12225 VN.n640 VN.n585 0.0389342
R12226 VN.n537 VN.n489 0.0389342
R12227 VN.n539 VN.n487 0.0389342
R12228 VN.n353 VN.n352 0.0338096
R12229 VN.n312 VN.n158 0.0338096
R12230 VN.n279 VN.n277 0.0338096
R12231 VN.n229 VN.n228 0.0338096
R12232 VN.n609 VN.n605 0.0338096
R12233 VN.n654 VN.n579 0.0338096
R12234 VN.n687 VN.n686 0.0338096
R12235 VN.n528 VN.n491 0.0338096
R12236 VN.n38 VN.n36 0.0325285
R12237 VN.n823 VN.n786 0.0325285
R12238 VN.n350 VN.n349 0.0325285
R12239 VN.n317 VN.n316 0.0325285
R12240 VN.n282 VN.n172 0.0325285
R12241 VN.n233 VN.n190 0.0325285
R12242 VN.n406 VN.n404 0.0325285
R12243 VN.n439 VN.n381 0.0325285
R12244 VN.n461 VN.n133 0.0325285
R12245 VN.n101 VN.n100 0.0325285
R12246 VN.n606 VN.n604 0.0325285
R12247 VN.n650 VN.n649 0.0325285
R12248 VN.n683 VN.n566 0.0325285
R12249 VN.n533 VN.n532 0.0325285
R12250 VN.n755 VN.n754 0.0325285
R12251 VN.n849 VN.n0 0.0325285
R12252 VN.n56 VN.n55 0.0318879
R12253 VN.n842 VN.n841 0.0318879
R12254 VN.n424 VN.n389 0.0318879
R12255 VN.n458 VN.n457 0.0318879
R12256 VN.n479 VN.n478 0.0318879
R12257 VN.n79 VN.n78 0.0318879
R12258 VN.n732 VN.n730 0.0318879
R12259 VN.n820 VN.n819 0.0318879
R12260 VN.n50 VN.n49 0.0312473
R12261 VN.n836 VN.n835 0.0312473
R12262 VN.n419 VN.n393 0.0312473
R12263 VN.n452 VN.n451 0.0312473
R12264 VN.n121 VN.n119 0.0312473
R12265 VN.n83 VN.n74 0.0312473
R12266 VN.n736 VN.n727 0.0312473
R12267 VN.n793 VN.n791 0.0312473
R12268 VN.n376 VN.n152 0.0306068
R12269 VN.n373 VN.n372 0.0306068
R12270 VN.n286 VN.n170 0.0306068
R12271 VN.n288 VN.n168 0.0306068
R12272 VN.n250 VN.n249 0.0306068
R12273 VN.n254 VN.n253 0.0306068
R12274 VN.n203 VN.n200 0.0306068
R12275 VN.n634 VN.n633 0.0306068
R12276 VN.n630 VN.n592 0.0306068
R12277 VN.n680 VN.n679 0.0306068
R12278 VN.n677 VN.n568 0.0306068
R12279 VN.n710 VN.n485 0.0306068
R12280 VN.n707 VN.n706 0.0306068
R12281 VN.n504 VN.n501 0.0306068
R12282 VN.n368 VN.n336 0.0299662
R12283 VN.n365 VN.n364 0.0299662
R12284 VN.n295 VN.n166 0.0299662
R12285 VN.n297 VN.n164 0.0299662
R12286 VN.n259 VN.n258 0.0299662
R12287 VN.n263 VN.n262 0.0299662
R12288 VN.n211 VN.n198 0.0299662
R12289 VN.n213 VN.n196 0.0299662
R12290 VN.n626 VN.n625 0.0299662
R12291 VN.n622 VN.n597 0.0299662
R12292 VN.n670 VN.n570 0.0299662
R12293 VN.n668 VN.n573 0.0299662
R12294 VN.n702 VN.n552 0.0299662
R12295 VN.n699 VN.n698 0.0299662
R12296 VN.n511 VN.n499 0.0299662
R12297 VN.n513 VN.n497 0.0299662
R12298 VN.n30 VN.n28 0.0270836
R12299 VN.n779 VN.n777 0.0270836
R12300 VN.n414 VN.n398 0.0270836
R12301 VN.n144 VN.n142 0.0270836
R12302 VN.n470 VN.n126 0.0270836
R12303 VN.n90 VN.n72 0.0270836
R12304 VN.n744 VN.n743 0.0270836
R12305 VN.n811 VN.n798 0.0270836
R12306 VN.n360 VN.n341 0.0258025
R12307 VN.n357 VN.n356 0.0258025
R12308 VN.n304 VN.n162 0.0258025
R12309 VN.n307 VN.n306 0.0258025
R12310 VN.n269 VN.n268 0.0258025
R12311 VN.n274 VN.n176 0.0258025
R12312 VN.n219 VN.n218 0.0258025
R12313 VN.n223 VN.n222 0.0258025
R12314 VN.n618 VN.n617 0.0258025
R12315 VN.n614 VN.n602 0.0258025
R12316 VN.n661 VN.n575 0.0258025
R12317 VN.n659 VN.n577 0.0258025
R12318 VN.n694 VN.n557 0.0258025
R12319 VN.n691 VN.n690 0.0258025
R12320 VN.n520 VN.n495 0.0258025
R12321 VN.n523 VN.n522 0.0258025
R12322 VN.n202 VN.n201 0.0170406
R12323 VN.n503 VN.n502 0.0170406
R12324 VN.n361 VN.n360 0.0149128
R12325 VN.n356 VN.n344 0.0149128
R12326 VN.n301 VN.n162 0.0149128
R12327 VN.n306 VN.n160 0.0149128
R12328 VN.n269 VN.n266 0.0149128
R12329 VN.n274 VN.n273 0.0149128
R12330 VN.n218 VN.n217 0.0149128
R12331 VN.n222 VN.n192 0.0149128
R12332 VN.n618 VN.n598 0.0149128
R12333 VN.n614 VN.n613 0.0149128
R12334 VN.n664 VN.n575 0.0149128
R12335 VN.n656 VN.n577 0.0149128
R12336 VN.n695 VN.n694 0.0149128
R12337 VN.n690 VN.n560 0.0149128
R12338 VN.n517 VN.n495 0.0149128
R12339 VN.n522 VN.n493 0.0149128
R12340 VN.n43 VN.n30 0.0136317
R12341 VN.n829 VN.n779 0.0136317
R12342 VN.n357 VN.n343 0.0136317
R12343 VN.n307 VN.n305 0.0136317
R12344 VN.n267 VN.n176 0.0136317
R12345 VN.n223 VN.n194 0.0136317
R12346 VN.n411 VN.n398 0.0136317
R12347 VN.n445 VN.n144 0.0136317
R12348 VN.n467 VN.n126 0.0136317
R12349 VN.n72 VN.n69 0.0136317
R12350 VN.n602 VN.n600 0.0136317
R12351 VN.n660 VN.n659 0.0136317
R12352 VN.n691 VN.n559 0.0136317
R12353 VN.n523 VN.n521 0.0136317
R12354 VN.n743 VN.n723 0.0136317
R12355 VN.n808 VN.n798 0.0136317
R12356 VN.n369 VN.n368 0.0107491
R12357 VN.n364 VN.n339 0.0107491
R12358 VN.n292 VN.n166 0.0107491
R12359 VN.n300 VN.n164 0.0107491
R12360 VN.n259 VN.n257 0.0107491
R12361 VN.n263 VN.n178 0.0107491
R12362 VN.n207 VN.n198 0.0107491
R12363 VN.n216 VN.n196 0.0107491
R12364 VN.n626 VN.n593 0.0107491
R12365 VN.n622 VN.n621 0.0107491
R12366 VN.n673 VN.n570 0.0107491
R12367 VN.n665 VN.n573 0.0107491
R12368 VN.n703 VN.n702 0.0107491
R12369 VN.n698 VN.n555 0.0107491
R12370 VN.n508 VN.n499 0.0107491
R12371 VN.n516 VN.n497 0.0107491
R12372 VN.n372 VN.n334 0.0101085
R12373 VN.n291 VN.n168 0.0101085
R12374 VN.n254 VN.n182 0.0101085
R12375 VN.n206 VN.n200 0.0101085
R12376 VN.n630 VN.n629 0.0101085
R12377 VN.n674 VN.n568 0.0101085
R12378 VN.n706 VN.n550 0.0101085
R12379 VN.n507 VN.n501 0.0101085
R12380 VN.n49 VN.n48 0.00946797
R12381 VN.n835 VN.n834 0.00946797
R12382 VN.n365 VN.n338 0.00946797
R12383 VN.n297 VN.n296 0.00946797
R12384 VN.n262 VN.n180 0.00946797
R12385 VN.n213 VN.n212 0.00946797
R12386 VN.n416 VN.n393 0.00946797
R12387 VN.n451 VN.n450 0.00946797
R12388 VN.n472 VN.n121 0.00946797
R12389 VN.n86 VN.n74 0.00946797
R12390 VN.n597 VN.n595 0.00946797
R12391 VN.n669 VN.n668 0.00946797
R12392 VN.n699 VN.n554 0.00946797
R12393 VN.n513 VN.n512 0.00946797
R12394 VN.n739 VN.n727 0.00946797
R12395 VN.n813 VN.n793 0.00946797
R12396 VN.n55 VN.n54 0.0088274
R12397 VN.n841 VN.n840 0.0088274
R12398 VN.n373 VN.n333 0.0088274
R12399 VN.n288 VN.n287 0.0088274
R12400 VN.n253 VN.n184 0.0088274
R12401 VN.n203 VN.n202 0.0088274
R12402 VN.n421 VN.n389 0.0088274
R12403 VN.n457 VN.n456 0.0088274
R12404 VN.n478 VN.n477 0.0088274
R12405 VN.n78 VN.n76 0.0088274
R12406 VN.n592 VN.n590 0.0088274
R12407 VN.n678 VN.n677 0.0088274
R12408 VN.n707 VN.n549 0.0088274
R12409 VN.n504 VN.n503 0.0088274
R12410 VN.n730 VN.n729 0.0088274
R12411 VN.n819 VN.n818 0.0088274
R12412 VN.n36 VN.n35 0.00818683
R12413 VN.n786 VN.n784 0.00818683
R12414 VN.n404 VN.n403 0.00818683
R12415 VN.n381 VN.n149 0.00818683
R12416 VN.n133 VN.n131 0.00818683
R12417 VN.n100 VN.n99 0.00818683
R12418 VN.n754 VN.n753 0.00818683
R12419 VN.n804 VN.n0 0.00818683
R12420 VN.n353 VN.n346 0.00690569
R12421 VN.n352 VN.n347 0.00690569
R12422 VN.n312 VN.n311 0.00690569
R12423 VN.n315 VN.n158 0.00690569
R12424 VN.n277 VN.n174 0.00690569
R12425 VN.n279 VN.n278 0.00690569
R12426 VN.n228 VN.n227 0.00690569
R12427 VN.n230 VN.n229 0.00690569
R12428 VN.n605 VN.n603 0.00690569
R12429 VN.n609 VN.n608 0.00690569
R12430 VN.n655 VN.n654 0.00690569
R12431 VN.n651 VN.n579 0.00690569
R12432 VN.n687 VN.n562 0.00690569
R12433 VN.n686 VN.n563 0.00690569
R12434 VN.n528 VN.n527 0.00690569
R12435 VN.n531 VN.n491 0.00690569
R12436 VN VN.n849 0.00306228
R12437 VN.n386 VN.n384 0.00185849
R12438 VN.n428 VN.n387 0.00185849
R12439 VN.n108 VN.n107 0.00185849
R12440 VN.n114 VN.n113 0.00185849
R12441 VN.n13 VN.n12 0.00185849
R12442 VN.n19 VN.n18 0.00185849
R12443 VN.n762 VN.n761 0.00185849
R12444 VN.n768 VN.n767 0.00185849
R12445 VN.n333 VN.n152 0.00178114
R12446 VN.n338 VN.n336 0.00178114
R12447 VN.n343 VN.n341 0.00178114
R12448 VN.n349 VN.n347 0.00178114
R12449 VN.n287 VN.n286 0.00178114
R12450 VN.n296 VN.n295 0.00178114
R12451 VN.n305 VN.n304 0.00178114
R12452 VN.n316 VN.n315 0.00178114
R12453 VN.n249 VN.n184 0.00178114
R12454 VN.n258 VN.n180 0.00178114
R12455 VN.n268 VN.n267 0.00178114
R12456 VN.n278 VN.n172 0.00178114
R12457 VN.n324 VN.n323 0.00178114
R12458 VN.n330 VN.n329 0.00178114
R12459 VN.n240 VN.n239 0.00178114
R12460 VN.n246 VN.n245 0.00178114
R12461 VN.n212 VN.n211 0.00178114
R12462 VN.n219 VN.n194 0.00178114
R12463 VN.n230 VN.n190 0.00178114
R12464 VN.n633 VN.n590 0.00178114
R12465 VN.n625 VN.n595 0.00178114
R12466 VN.n617 VN.n600 0.00178114
R12467 VN.n608 VN.n606 0.00178114
R12468 VN.n679 VN.n678 0.00178114
R12469 VN.n670 VN.n669 0.00178114
R12470 VN.n661 VN.n660 0.00178114
R12471 VN.n651 VN.n650 0.00178114
R12472 VN.n549 VN.n485 0.00178114
R12473 VN.n554 VN.n552 0.00178114
R12474 VN.n559 VN.n557 0.00178114
R12475 VN.n566 VN.n563 0.00178114
R12476 VN.n585 VN.n583 0.00178114
R12477 VN.n638 VN.n586 0.00178114
R12478 VN.n540 VN.n539 0.00178114
R12479 VN.n546 VN.n545 0.00178114
R12480 VN.n512 VN.n511 0.00178114
R12481 VN.n521 VN.n520 0.00178114
R12482 VN.n532 VN.n531 0.00178114
R12483 a_n13990_n5465.n168 a_n13990_n5465.n167 9.23995
R12484 a_n13990_n5465.n31 a_n13990_n5465.n27 7.94229
R12485 a_n13990_n5465.n210 a_n13990_n5465.n207 7.94229
R12486 a_n13990_n5465.n166 a_n13990_n5465.t32 6.72766
R12487 a_n13990_n5465.n139 a_n13990_n5465.n134 6.58329
R12488 a_n13990_n5465.n174 a_n13990_n5465.n168 6.01251
R12489 a_n13990_n5465.n138 a_n13990_n5465.n137 5.85326
R12490 a_n13990_n5465.n131 a_n13990_n5465.n130 5.85326
R12491 a_n13990_n5465.n138 a_n13990_n5465.n136 5.84661
R12492 a_n13990_n5465.n26 a_n13990_n5465.n25 5.69423
R12493 a_n13990_n5465.n33 a_n13990_n5465.n32 5.69423
R12494 a_n13990_n5465.n206 a_n13990_n5465.n205 5.69423
R12495 a_n13990_n5465.n212 a_n13990_n5465.n211 5.69423
R12496 a_n13990_n5465.n26 a_n13990_n5465.n24 5.49558
R12497 a_n13990_n5465.n206 a_n13990_n5465.n204 5.49558
R12498 a_n13990_n5465.n0 a_n13990_n5465.n218 4.22068
R12499 a_n13990_n5465.t51 a_n13990_n5465.n1 5.69068
R12500 a_n13990_n5465.n216 a_n13990_n5465.n2 4.22068
R12501 a_n13990_n5465.n3 a_n13990_n5465.n172 4.22068
R12502 a_n13990_n5465.t69 a_n13990_n5465.n4 5.69068
R12503 a_n13990_n5465.n170 a_n13990_n5465.n5 4.22068
R12504 a_n13990_n5465.n7 a_n13990_n5465.n88 4.58971
R12505 a_n13990_n5465.n8 a_n13990_n5465.t11 5.84971
R12506 a_n13990_n5465.n9 a_n13990_n5465.n96 4.58971
R12507 a_n13990_n5465.n6 a_n13990_n5465.n142 5.47076
R12508 a_n13990_n5465.n134 a_n13990_n5465.n133 4.59326
R12509 a_n13990_n5465.n167 a_n13990_n5465.n166 4.52463
R12510 a_n13990_n5465.n146 a_n13990_n5465.t34 4.41563
R12511 a_n13990_n5465.n161 a_n13990_n5465.n159 4.41563
R12512 a_n13990_n5465.n31 a_n13990_n5465.n30 4.22423
R12513 a_n13990_n5465.n210 a_n13990_n5465.n209 4.22423
R12514 a_n13990_n5465.n166 a_n13990_n5465.n165 4.21432
R12515 a_n13990_n5465.n124 a_n13990_n5465.n123 4.21195
R12516 a_n13990_n5465.n126 a_n13990_n5465.t22 4.21195
R12517 a_n13990_n5465.n103 a_n13990_n5465.n102 4.21195
R12518 a_n13990_n5465.n99 a_n13990_n5465.t0 4.21195
R12519 a_n13990_n5465.n10 a_n13990_n5465.t120 4.05054
R12520 a_n13990_n5465.n223 a_n13990_n5465.t81 4.05054
R12521 a_n13990_n5465.n45 a_n13990_n5465.n44 4.05054
R12522 a_n13990_n5465.n47 a_n13990_n5465.t70 4.05054
R12523 a_n13990_n5465.n57 a_n13990_n5465.n56 4.05054
R12524 a_n13990_n5465.n59 a_n13990_n5465.t113 4.05054
R12525 a_n13990_n5465.n36 a_n13990_n5465.n35 4.05054
R12526 a_n13990_n5465.n73 a_n13990_n5465.t121 4.05054
R12527 a_n13990_n5465.n82 a_n13990_n5465.n81 4.05054
R12528 a_n13990_n5465.n84 a_n13990_n5465.t105 4.05054
R12529 a_n13990_n5465.n185 a_n13990_n5465.n184 4.05054
R12530 a_n13990_n5465.n187 a_n13990_n5465.t66 4.05054
R12531 a_n13990_n5465.n197 a_n13990_n5465.n196 4.05054
R12532 a_n13990_n5465.n199 a_n13990_n5465.t88 4.05054
R12533 a_n13990_n5465.n66 a_n13990_n5465.n65 4.05054
R12534 a_n13990_n5465.n228 a_n13990_n5465.n227 4.05054
R12535 a_n13990_n5465.n124 a_n13990_n5465.n122 4.03668
R12536 a_n13990_n5465.n126 a_n13990_n5465.t139 4.03668
R12537 a_n13990_n5465.n103 a_n13990_n5465.n101 4.03668
R12538 a_n13990_n5465.n99 a_n13990_n5465.t5 4.03668
R12539 a_n13990_n5465.n227 a_n13990_n5465.n226 3.87765
R12540 a_n13990_n5465.n10 a_n13990_n5465.t119 3.87765
R12541 a_n13990_n5465.n223 a_n13990_n5465.t79 3.87765
R12542 a_n13990_n5465.n45 a_n13990_n5465.n43 3.87765
R12543 a_n13990_n5465.n47 a_n13990_n5465.t67 3.87765
R12544 a_n13990_n5465.n57 a_n13990_n5465.n55 3.87765
R12545 a_n13990_n5465.n59 a_n13990_n5465.t112 3.87765
R12546 a_n13990_n5465.n36 a_n13990_n5465.n34 3.87765
R12547 a_n13990_n5465.n73 a_n13990_n5465.t124 3.87765
R12548 a_n13990_n5465.n82 a_n13990_n5465.n80 3.87765
R12549 a_n13990_n5465.n84 a_n13990_n5465.t107 3.87765
R12550 a_n13990_n5465.n185 a_n13990_n5465.n183 3.87765
R12551 a_n13990_n5465.n187 a_n13990_n5465.t68 3.87765
R12552 a_n13990_n5465.n197 a_n13990_n5465.n195 3.87765
R12553 a_n13990_n5465.n199 a_n13990_n5465.t89 3.87765
R12554 a_n13990_n5465.n66 a_n13990_n5465.n64 3.87765
R12555 a_n13990_n5465.n146 a_n13990_n5465.t30 3.833
R12556 a_n13990_n5465.n161 a_n13990_n5465.n160 3.833
R12557 a_n13990_n5465.n116 a_n13990_n5465.n110 3.81703
R12558 a_n13990_n5465.n97 a_n13990_n5465.n9 3.95161
R12559 a_n13990_n5465.n158 a_n13990_n5465.n152 3.80578
R12560 a_n13990_n5465.n145 a_n13990_n5465.n6 3.90344
R12561 a_n13990_n5465.n141 a_n13990_n5465.n140 3.69568
R12562 a_n13990_n5465.n62 a_n13990_n5465.n33 3.25667
R12563 a_n13990_n5465.n151 a_n13990_n5465.n148 3.15563
R12564 a_n13990_n5465.n157 a_n13990_n5465.n154 3.15563
R12565 a_n13990_n5465.n2 a_n13990_n5465.n214 3.15553
R12566 a_n13990_n5465.n5 a_n13990_n5465.n63 3.15553
R12567 a_n13990_n5465.n121 a_n13990_n5465.n120 2.95195
R12568 a_n13990_n5465.n115 a_n13990_n5465.n114 2.95195
R12569 a_n13990_n5465.n109 a_n13990_n5465.n108 2.95195
R12570 a_n13990_n5465.n94 a_n13990_n5465.n93 2.95195
R12571 a_n13990_n5465.n121 a_n13990_n5465.n118 2.77668
R12572 a_n13990_n5465.n115 a_n13990_n5465.n112 2.77668
R12573 a_n13990_n5465.n109 a_n13990_n5465.n106 2.77668
R12574 a_n13990_n5465.n94 a_n13990_n5465.n91 2.77668
R12575 a_n13990_n5465.n72 a_n13990_n5465.n66 2.73714
R12576 a_n13990_n5465.n42 a_n13990_n5465.n36 2.73714
R12577 a_n13990_n5465.n16 a_n13990_n5465.n10 2.73672
R12578 a_n13990_n5465.n79 a_n13990_n5465.n73 2.73672
R12579 a_n13990_n5465.n152 a_n13990_n5465.n146 2.71872
R12580 a_n13990_n5465.n125 a_n13990_n5465.n121 2.71872
R12581 a_n13990_n5465.n188 a_n13990_n5465.n186 2.60203
R12582 a_n13990_n5465.n48 a_n13990_n5465.n46 2.60203
R12583 a_n13990_n5465.n141 a_n13990_n5465.n86 2.5825
R12584 a_n13990_n5465.n15 a_n13990_n5465.n14 2.58054
R12585 a_n13990_n5465.n21 a_n13990_n5465.n20 2.58054
R12586 a_n13990_n5465.n53 a_n13990_n5465.n52 2.58054
R12587 a_n13990_n5465.n41 a_n13990_n5465.n40 2.58054
R12588 a_n13990_n5465.n78 a_n13990_n5465.n77 2.58054
R12589 a_n13990_n5465.n181 a_n13990_n5465.n180 2.58054
R12590 a_n13990_n5465.n193 a_n13990_n5465.n192 2.58054
R12591 a_n13990_n5465.n71 a_n13990_n5465.n70 2.58054
R12592 a_n13990_n5465.n151 a_n13990_n5465.n150 2.573
R12593 a_n13990_n5465.n157 a_n13990_n5465.n156 2.573
R12594 a_n13990_n5465.n104 a_n13990_n5465.n100 2.56118
R12595 a_n13990_n5465.n127 a_n13990_n5465.n125 2.56118
R12596 a_n13990_n5465.n131 a_n13990_n5465.n86 2.54573
R12597 a_n13990_n5465.n200 a_n13990_n5465.n198 2.53418
R12598 a_n13990_n5465.n85 a_n13990_n5465.n83 2.53418
R12599 a_n13990_n5465.n60 a_n13990_n5465.n58 2.53418
R12600 a_n13990_n5465.n225 a_n13990_n5465.n224 2.53418
R12601 a_n13990_n5465.n213 a_n13990_n5465.n212 2.51873
R12602 a_n13990_n5465.n15 a_n13990_n5465.n12 2.40765
R12603 a_n13990_n5465.n21 a_n13990_n5465.n18 2.40765
R12604 a_n13990_n5465.n53 a_n13990_n5465.n50 2.40765
R12605 a_n13990_n5465.n41 a_n13990_n5465.n38 2.40765
R12606 a_n13990_n5465.n78 a_n13990_n5465.n75 2.40765
R12607 a_n13990_n5465.n181 a_n13990_n5465.n178 2.40765
R12608 a_n13990_n5465.n193 a_n13990_n5465.n190 2.40765
R12609 a_n13990_n5465.n71 a_n13990_n5465.n68 2.40765
R12610 a_n13990_n5465.n129 a_n13990_n5465.n89 2.27857
R12611 a_n13990_n5465.n221 a_n13990_n5465.n27 2.23844
R12612 a_n13990_n5465.n98 a_n13990_n5465.n94 2.00466
R12613 a_n13990_n5465.n163 a_n13990_n5465.n162 1.67718
R12614 a_n13990_n5465.n89 a_n13990_n5465.n7 1.67353
R12615 a_n13990_n5465.n219 a_n13990_n5465.n0 1.65553
R12616 a_n13990_n5465.n173 a_n13990_n5465.n3 1.65553
R12617 a_n13990_n5465.n202 a_n13990_n5465.n201 1.5005
R12618 a_n13990_n5465.n98 a_n13990_n5465.n97 1.5005
R12619 a_n13990_n5465.n129 a_n13990_n5465.n128 1.5005
R12620 a_n13990_n5465.n140 a_n13990_n5465.n139 1.5005
R12621 a_n13990_n5465.n174 a_n13990_n5465.n173 1.5005
R12622 a_n13990_n5465.n176 a_n13990_n5465.n175 1.5005
R12623 a_n13990_n5465.n207 a_n13990_n5465.n28 1.5005
R12624 a_n13990_n5465.n220 a_n13990_n5465.n219 1.5005
R12625 a_n13990_n5465.n222 a_n13990_n5465.n221 1.5005
R12626 a_n13990_n5465.n62 a_n13990_n5465.n61 1.5005
R12627 a_n13990_n5465.n12 a_n13990_n5465.t48 1.4705
R12628 a_n13990_n5465.n12 a_n13990_n5465.n11 1.4705
R12629 a_n13990_n5465.n14 a_n13990_n5465.t50 1.4705
R12630 a_n13990_n5465.n14 a_n13990_n5465.n13 1.4705
R12631 a_n13990_n5465.n18 a_n13990_n5465.t122 1.4705
R12632 a_n13990_n5465.n18 a_n13990_n5465.n17 1.4705
R12633 a_n13990_n5465.n20 a_n13990_n5465.t126 1.4705
R12634 a_n13990_n5465.n20 a_n13990_n5465.n19 1.4705
R12635 a_n13990_n5465.n50 a_n13990_n5465.t104 1.4705
R12636 a_n13990_n5465.n50 a_n13990_n5465.n49 1.4705
R12637 a_n13990_n5465.n52 a_n13990_n5465.t106 1.4705
R12638 a_n13990_n5465.n52 a_n13990_n5465.n51 1.4705
R12639 a_n13990_n5465.n38 a_n13990_n5465.t63 1.4705
R12640 a_n13990_n5465.n38 a_n13990_n5465.n37 1.4705
R12641 a_n13990_n5465.n40 a_n13990_n5465.t65 1.4705
R12642 a_n13990_n5465.n40 a_n13990_n5465.n39 1.4705
R12643 a_n13990_n5465.n24 a_n13990_n5465.t53 1.4705
R12644 a_n13990_n5465.n24 a_n13990_n5465.n23 1.4705
R12645 a_n13990_n5465.n30 a_n13990_n5465.t91 1.4705
R12646 a_n13990_n5465.n30 a_n13990_n5465.n29 1.4705
R12647 a_n13990_n5465.n218 a_n13990_n5465.t90 1.4705
R12648 a_n13990_n5465.n218 a_n13990_n5465.n217 1.4705
R12649 a_n13990_n5465.n216 a_n13990_n5465.t49 1.4705
R12650 a_n13990_n5465.n216 a_n13990_n5465.n215 1.4705
R12651 a_n13990_n5465.n204 a_n13990_n5465.t80 1.4705
R12652 a_n13990_n5465.n204 a_n13990_n5465.n203 1.4705
R12653 a_n13990_n5465.n209 a_n13990_n5465.t108 1.4705
R12654 a_n13990_n5465.n209 a_n13990_n5465.n208 1.4705
R12655 a_n13990_n5465.n75 a_n13990_n5465.t72 1.4705
R12656 a_n13990_n5465.n75 a_n13990_n5465.n74 1.4705
R12657 a_n13990_n5465.n77 a_n13990_n5465.t71 1.4705
R12658 a_n13990_n5465.n77 a_n13990_n5465.n76 1.4705
R12659 a_n13990_n5465.n178 a_n13990_n5465.t118 1.4705
R12660 a_n13990_n5465.n178 a_n13990_n5465.n177 1.4705
R12661 a_n13990_n5465.n180 a_n13990_n5465.t117 1.4705
R12662 a_n13990_n5465.n180 a_n13990_n5465.n179 1.4705
R12663 a_n13990_n5465.n190 a_n13990_n5465.t76 1.4705
R12664 a_n13990_n5465.n190 a_n13990_n5465.n189 1.4705
R12665 a_n13990_n5465.n192 a_n13990_n5465.t75 1.4705
R12666 a_n13990_n5465.n192 a_n13990_n5465.n191 1.4705
R12667 a_n13990_n5465.n68 a_n13990_n5465.t111 1.4705
R12668 a_n13990_n5465.n68 a_n13990_n5465.n67 1.4705
R12669 a_n13990_n5465.n70 a_n13990_n5465.t110 1.4705
R12670 a_n13990_n5465.n70 a_n13990_n5465.n69 1.4705
R12671 a_n13990_n5465.n172 a_n13990_n5465.t98 1.4705
R12672 a_n13990_n5465.n172 a_n13990_n5465.n171 1.4705
R12673 a_n13990_n5465.n170 a_n13990_n5465.t101 1.4705
R12674 a_n13990_n5465.n170 a_n13990_n5465.n169 1.4705
R12675 a_n13990_n5465.n16 a_n13990_n5465.n15 1.46537
R12676 a_n13990_n5465.n227 a_n13990_n5465.n225 1.46537
R12677 a_n13990_n5465.n22 a_n13990_n5465.n21 1.46537
R12678 a_n13990_n5465.n46 a_n13990_n5465.n45 1.46537
R12679 a_n13990_n5465.n48 a_n13990_n5465.n47 1.46537
R12680 a_n13990_n5465.n54 a_n13990_n5465.n53 1.46537
R12681 a_n13990_n5465.n58 a_n13990_n5465.n57 1.46537
R12682 a_n13990_n5465.n42 a_n13990_n5465.n41 1.46537
R12683 a_n13990_n5465.n79 a_n13990_n5465.n78 1.46537
R12684 a_n13990_n5465.n83 a_n13990_n5465.n82 1.46537
R12685 a_n13990_n5465.n182 a_n13990_n5465.n181 1.46537
R12686 a_n13990_n5465.n186 a_n13990_n5465.n185 1.46537
R12687 a_n13990_n5465.n188 a_n13990_n5465.n187 1.46537
R12688 a_n13990_n5465.n194 a_n13990_n5465.n193 1.46537
R12689 a_n13990_n5465.n198 a_n13990_n5465.n197 1.46537
R12690 a_n13990_n5465.n72 a_n13990_n5465.n71 1.46537
R12691 a_n13990_n5465.n125 a_n13990_n5465.n124 1.46537
R12692 a_n13990_n5465.n116 a_n13990_n5465.n115 1.46537
R12693 a_n13990_n5465.n110 a_n13990_n5465.n109 1.46537
R12694 a_n13990_n5465.n104 a_n13990_n5465.n103 1.46537
R12695 a_n13990_n5465.n152 a_n13990_n5465.n151 1.46537
R12696 a_n13990_n5465.n158 a_n13990_n5465.n157 1.46537
R12697 a_n13990_n5465.n162 a_n13990_n5465.n161 1.46537
R12698 a_n13990_n5465.n224 a_n13990_n5465.n223 1.46535
R12699 a_n13990_n5465.n60 a_n13990_n5465.n59 1.46535
R12700 a_n13990_n5465.n85 a_n13990_n5465.n84 1.46535
R12701 a_n13990_n5465.n200 a_n13990_n5465.n199 1.46535
R12702 a_n13990_n5465.n127 a_n13990_n5465.n126 1.46535
R12703 a_n13990_n5465.n100 a_n13990_n5465.n99 1.46535
R12704 a_n13990_n5465.n168 a_n13990_n5465.n63 1.43535
R12705 a_n13990_n5465.n145 a_n13990_n5465.n141 1.31908
R12706 a_n13990_n5465.n225 a_n13990_n5465.n16 1.27228
R12707 a_n13990_n5465.n33 a_n13990_n5465.n31 1.27228
R12708 a_n13990_n5465.n212 a_n13990_n5465.n210 1.27228
R12709 a_n13990_n5465.n198 a_n13990_n5465.n194 1.27228
R12710 a_n13990_n5465.n194 a_n13990_n5465.n188 1.27228
R12711 a_n13990_n5465.n186 a_n13990_n5465.n182 1.27228
R12712 a_n13990_n5465.n83 a_n13990_n5465.n79 1.27228
R12713 a_n13990_n5465.n58 a_n13990_n5465.n54 1.27228
R12714 a_n13990_n5465.n54 a_n13990_n5465.n48 1.27228
R12715 a_n13990_n5465.n46 a_n13990_n5465.n22 1.27228
R12716 a_n13990_n5465.n148 a_n13990_n5465.t35 1.2605
R12717 a_n13990_n5465.n148 a_n13990_n5465.n147 1.2605
R12718 a_n13990_n5465.n150 a_n13990_n5465.t31 1.2605
R12719 a_n13990_n5465.n150 a_n13990_n5465.n149 1.2605
R12720 a_n13990_n5465.n154 a_n13990_n5465.t28 1.2605
R12721 a_n13990_n5465.n154 a_n13990_n5465.n153 1.2605
R12722 a_n13990_n5465.n156 a_n13990_n5465.t36 1.2605
R12723 a_n13990_n5465.n156 a_n13990_n5465.n155 1.2605
R12724 a_n13990_n5465.n165 a_n13990_n5465.t33 1.2605
R12725 a_n13990_n5465.n165 a_n13990_n5465.n164 1.2605
R12726 a_n13990_n5465.n144 a_n13990_n5465.t29 1.2605
R12727 a_n13990_n5465.n144 a_n13990_n5465.n143 1.2605
R12728 a_n13990_n5465.n88 a_n13990_n5465.t15 1.2605
R12729 a_n13990_n5465.n88 a_n13990_n5465.n87 1.2605
R12730 a_n13990_n5465.n96 a_n13990_n5465.t10 1.2605
R12731 a_n13990_n5465.n96 a_n13990_n5465.n95 1.2605
R12732 a_n13990_n5465.n136 a_n13990_n5465.t8 1.2605
R12733 a_n13990_n5465.n136 a_n13990_n5465.n135 1.2605
R12734 a_n13990_n5465.n133 a_n13990_n5465.t17 1.2605
R12735 a_n13990_n5465.n133 a_n13990_n5465.n132 1.2605
R12736 a_n13990_n5465.n118 a_n13990_n5465.t7 1.2605
R12737 a_n13990_n5465.n118 a_n13990_n5465.n117 1.2605
R12738 a_n13990_n5465.n120 a_n13990_n5465.t20 1.2605
R12739 a_n13990_n5465.n120 a_n13990_n5465.n119 1.2605
R12740 a_n13990_n5465.n112 a_n13990_n5465.t1 1.2605
R12741 a_n13990_n5465.n112 a_n13990_n5465.n111 1.2605
R12742 a_n13990_n5465.n114 a_n13990_n5465.t24 1.2605
R12743 a_n13990_n5465.n114 a_n13990_n5465.n113 1.2605
R12744 a_n13990_n5465.n106 a_n13990_n5465.t21 1.2605
R12745 a_n13990_n5465.n106 a_n13990_n5465.n105 1.2605
R12746 a_n13990_n5465.n108 a_n13990_n5465.t4 1.2605
R12747 a_n13990_n5465.n108 a_n13990_n5465.n107 1.2605
R12748 a_n13990_n5465.n91 a_n13990_n5465.t27 1.2605
R12749 a_n13990_n5465.n91 a_n13990_n5465.n90 1.2605
R12750 a_n13990_n5465.n93 a_n13990_n5465.t25 1.2605
R12751 a_n13990_n5465.n93 a_n13990_n5465.n92 1.2605
R12752 a_n13990_n5465.n134 a_n13990_n5465.n131 1.25428
R12753 a_n13990_n5465.n110 a_n13990_n5465.n104 1.25428
R12754 a_n13990_n5465.n162 a_n13990_n5465.n158 1.25428
R12755 a_n13990_n5465.n139 a_n13990_n5465.n138 1.04573
R12756 a_n13990_n5465.n27 a_n13990_n5465.n26 1.01873
R12757 a_n13990_n5465.n207 a_n13990_n5465.n206 1.01873
R12758 a_n13990_n5465.n214 a_n13990_n5465.n62 0.778574
R12759 a_n13990_n5465.n202 a_n13990_n5465.n63 0.778574
R12760 a_n13990_n5465.n221 a_n13990_n5465.n220 0.778574
R12761 a_n13990_n5465.n175 a_n13990_n5465.n174 0.778574
R12762 a_n13990_n5465.n213 a_n13990_n5465.n202 0.738439
R12763 a_n13990_n5465.n97 a_n13990_n5465.n86 0.738439
R12764 a_n13990_n5465.n140 a_n13990_n5465.n129 0.738439
R12765 a_n13990_n5465.n175 a_n13990_n5465.n28 0.738439
R12766 a_n13990_n5465.n167 a_n13990_n5465.n163 0.737223
R12767 a_n13990_n5465.n201 a_n13990_n5465.n200 0.699581
R12768 a_n13990_n5465.n176 a_n13990_n5465.n85 0.699581
R12769 a_n13990_n5465.n100 a_n13990_n5465.n98 0.699581
R12770 a_n13990_n5465.n128 a_n13990_n5465.n127 0.699581
R12771 a_n13990_n5465.n61 a_n13990_n5465.n60 0.699581
R12772 a_n13990_n5465.n224 a_n13990_n5465.n222 0.699581
R12773 a_n13990_n5465.n163 a_n13990_n5465.n145 0.585196
R12774 a_n13990_n5465.n201 a_n13990_n5465.n72 0.557791
R12775 a_n13990_n5465.n182 a_n13990_n5465.n176 0.557791
R12776 a_n13990_n5465.n61 a_n13990_n5465.n42 0.557791
R12777 a_n13990_n5465.n222 a_n13990_n5465.n22 0.557791
R12778 a_n13990_n5465.n128 a_n13990_n5465.n116 0.539791
R12779 a_n13990_n5465.n214 a_n13990_n5465.n213 0.530466
R12780 a_n13990_n5465.n220 a_n13990_n5465.n28 0.530466
R12781 a_n13990_n5465.n1 a_n13990_n5465.n2 1.27228
R12782 a_n13990_n5465.n219 a_n13990_n5465.n1 7.30549
R12783 a_n13990_n5465.t85 a_n13990_n5465.n0 6.96214
R12784 a_n13990_n5465.n4 a_n13990_n5465.n5 1.27228
R12785 a_n13990_n5465.n173 a_n13990_n5465.n4 7.30549
R12786 a_n13990_n5465.t125 a_n13990_n5465.n3 6.96214
R12787 a_n13990_n5465.n144 a_n13990_n5465.n6 5.45652
R12788 a_n13990_n5465.n8 a_n13990_n5465.n9 1.25428
R12789 a_n13990_n5465.n89 a_n13990_n5465.n8 5.95549
R12790 a_n13990_n5465.t16 a_n13990_n5465.n7 7.10317
R12791 a_5396_9163.n45 a_5396_9163.n40 7.94229
R12792 a_5396_9163.n105 a_5396_9163.n102 7.94229
R12793 a_5396_9163.n141 a_5396_9163.t107 6.58663
R12794 a_5396_9163.n202 a_5396_9163.t102 6.58663
R12795 a_5396_9163.n269 a_5396_9163.n268 5.95439
R12796 a_5396_9163.n204 a_5396_9163.n203 5.95439
R12797 a_5396_9163.n44 a_5396_9163.n43 5.69423
R12798 a_5396_9163.n37 a_5396_9163.n36 5.69423
R12799 a_5396_9163.n101 a_5396_9163.n100 5.69423
R12800 a_5396_9163.n107 a_5396_9163.n106 5.69423
R12801 a_5396_9163.n44 a_5396_9163.n42 5.49558
R12802 a_5396_9163.n101 a_5396_9163.n99 5.49558
R12803 a_5396_9163.n269 a_5396_9163.t90 5.31528
R12804 a_5396_9163.n204 a_5396_9163.t110 5.31528
R12805 a_5396_9163.n0 a_5396_9163.n35 4.22068
R12806 a_5396_9163.n1 a_5396_9163.t82 5.69068
R12807 a_5396_9163.n2 a_5396_9163.n33 4.22068
R12808 a_5396_9163.n3 a_5396_9163.n279 4.22068
R12809 a_5396_9163.t13 a_5396_9163.n4 5.69068
R12810 a_5396_9163.n277 a_5396_9163.n5 4.22068
R12811 a_5396_9163.n168 a_5396_9163.n7 3.84173
R12812 a_5396_9163.n212 a_5396_9163.n10 3.84173
R12813 a_5396_9163.n6 a_5396_9163.n169 5.31173
R12814 a_5396_9163.n166 a_5396_9163.n8 5.31173
R12815 a_5396_9163.n9 a_5396_9163.n213 5.31173
R12816 a_5396_9163.n210 a_5396_9163.n11 5.31173
R12817 a_5396_9163.n273 a_5396_9163.n272 4.50663
R12818 a_5396_9163.n208 a_5396_9163.n207 4.50663
R12819 a_5396_9163.n199 a_5396_9163.n8 4.46113
R12820 a_5396_9163.n40 a_5396_9163.n39 4.22423
R12821 a_5396_9163.n105 a_5396_9163.n104 4.22423
R12822 a_5396_9163.n12 a_5396_9163.t84 4.05054
R12823 a_5396_9163.n21 a_5396_9163.n20 4.05054
R12824 a_5396_9163.n120 a_5396_9163.n119 4.05054
R12825 a_5396_9163.n122 a_5396_9163.t46 4.05054
R12826 a_5396_9163.n132 a_5396_9163.n131 4.05054
R12827 a_5396_9163.n134 a_5396_9163.t52 4.05054
R12828 a_5396_9163.n111 a_5396_9163.n110 4.05054
R12829 a_5396_9163.n80 a_5396_9163.t42 4.05054
R12830 a_5396_9163.n89 a_5396_9163.n88 4.05054
R12831 a_5396_9163.n91 a_5396_9163.t18 4.05054
R12832 a_5396_9163.n72 a_5396_9163.n71 4.05054
R12833 a_5396_9163.n68 a_5396_9163.t54 4.05054
R12834 a_5396_9163.n60 a_5396_9163.n59 4.05054
R12835 a_5396_9163.n56 a_5396_9163.t28 4.05054
R12836 a_5396_9163.n48 a_5396_9163.n47 4.05054
R12837 a_5396_9163.t87 a_5396_9163.n285 4.05054
R12838 a_5396_9163.n274 a_5396_9163.n30 3.97558
R12839 a_5396_9163.n285 a_5396_9163.t50 3.87765
R12840 a_5396_9163.n12 a_5396_9163.t73 3.87765
R12841 a_5396_9163.n21 a_5396_9163.n19 3.87765
R12842 a_5396_9163.n120 a_5396_9163.n118 3.87765
R12843 a_5396_9163.n122 a_5396_9163.t83 3.87765
R12844 a_5396_9163.n132 a_5396_9163.n130 3.87765
R12845 a_5396_9163.n134 a_5396_9163.t59 3.87765
R12846 a_5396_9163.n111 a_5396_9163.n109 3.87765
R12847 a_5396_9163.n80 a_5396_9163.t35 3.87765
R12848 a_5396_9163.n89 a_5396_9163.n87 3.87765
R12849 a_5396_9163.n91 a_5396_9163.t10 3.87765
R12850 a_5396_9163.n72 a_5396_9163.n70 3.87765
R12851 a_5396_9163.n68 a_5396_9163.t49 3.87765
R12852 a_5396_9163.n60 a_5396_9163.n58 3.87765
R12853 a_5396_9163.n56 a_5396_9163.t22 3.87765
R12854 a_5396_9163.n48 a_5396_9163.n46 3.87765
R12855 a_5396_9163.n141 a_5396_9163.n140 3.84528
R12856 a_5396_9163.n272 a_5396_9163.n271 3.84528
R12857 a_5396_9163.n202 a_5396_9163.n201 3.84528
R12858 a_5396_9163.n207 a_5396_9163.n206 3.84528
R12859 a_5396_9163.n235 a_5396_9163.n229 3.79678
R12860 a_5396_9163.n258 a_5396_9163.n252 3.79678
R12861 a_5396_9163.n192 a_5396_9163.n186 3.79678
R12862 a_5396_9163.n159 a_5396_9163.n153 3.79678
R12863 a_5396_9163.n11 a_5396_9163.n209 3.87644
R12864 a_5396_9163.n265 a_5396_9163.n241 3.73034
R12865 a_5396_9163.n180 a_5396_9163.n174 3.73034
R12866 a_5396_9163.n37 a_5396_9163.n31 3.25667
R12867 a_5396_9163.n97 a_5396_9163.n2 3.15553
R12868 a_5396_9163.n5 a_5396_9163.n275 3.15553
R12869 a_5396_9163.n268 a_5396_9163.n141 3.00663
R12870 a_5396_9163.n203 a_5396_9163.n202 3.00663
R12871 a_5396_9163.n246 a_5396_9163.n243 2.7866
R12872 a_5396_9163.n251 a_5396_9163.n248 2.7866
R12873 a_5396_9163.n257 a_5396_9163.n254 2.7866
R12874 a_5396_9163.n263 a_5396_9163.n260 2.7866
R12875 a_5396_9163.n240 a_5396_9163.n237 2.7866
R12876 a_5396_9163.n234 a_5396_9163.n231 2.7866
R12877 a_5396_9163.n228 a_5396_9163.n225 2.7866
R12878 a_5396_9163.n222 a_5396_9163.n219 2.7866
R12879 a_5396_9163.n147 a_5396_9163.n144 2.7866
R12880 a_5396_9163.n152 a_5396_9163.n149 2.7866
R12881 a_5396_9163.n158 a_5396_9163.n155 2.7866
R12882 a_5396_9163.n164 a_5396_9163.n161 2.7866
R12883 a_5396_9163.n179 a_5396_9163.n176 2.7866
R12884 a_5396_9163.n185 a_5396_9163.n182 2.7866
R12885 a_5396_9163.n191 a_5396_9163.n188 2.7866
R12886 a_5396_9163.n197 a_5396_9163.n194 2.7866
R12887 a_5396_9163.n54 a_5396_9163.n48 2.73714
R12888 a_5396_9163.n117 a_5396_9163.n111 2.73714
R12889 a_5396_9163.n18 a_5396_9163.n12 2.73672
R12890 a_5396_9163.n86 a_5396_9163.n80 2.73672
R12891 a_5396_9163.n252 a_5396_9163.n246 2.73672
R12892 a_5396_9163.n153 a_5396_9163.n147 2.73672
R12893 a_5396_9163.n73 a_5396_9163.n69 2.60203
R12894 a_5396_9163.n123 a_5396_9163.n121 2.60203
R12895 a_5396_9163.n17 a_5396_9163.n16 2.58054
R12896 a_5396_9163.n27 a_5396_9163.n26 2.58054
R12897 a_5396_9163.n128 a_5396_9163.n127 2.58054
R12898 a_5396_9163.n116 a_5396_9163.n115 2.58054
R12899 a_5396_9163.n85 a_5396_9163.n84 2.58054
R12900 a_5396_9163.n78 a_5396_9163.n77 2.58054
R12901 a_5396_9163.n66 a_5396_9163.n65 2.58054
R12902 a_5396_9163.n53 a_5396_9163.n52 2.58054
R12903 a_5396_9163.n284 a_5396_9163.n22 2.53418
R12904 a_5396_9163.n61 a_5396_9163.n57 2.53418
R12905 a_5396_9163.n92 a_5396_9163.n90 2.53418
R12906 a_5396_9163.n135 a_5396_9163.n133 2.53418
R12907 a_5396_9163.n108 a_5396_9163.n107 2.51873
R12908 a_5396_9163.n17 a_5396_9163.n14 2.40765
R12909 a_5396_9163.n27 a_5396_9163.n24 2.40765
R12910 a_5396_9163.n128 a_5396_9163.n125 2.40765
R12911 a_5396_9163.n116 a_5396_9163.n113 2.40765
R12912 a_5396_9163.n85 a_5396_9163.n82 2.40765
R12913 a_5396_9163.n78 a_5396_9163.n75 2.40765
R12914 a_5396_9163.n66 a_5396_9163.n63 2.40765
R12915 a_5396_9163.n53 a_5396_9163.n50 2.40765
R12916 a_5396_9163.n216 a_5396_9163.n9 2.37644
R12917 a_5396_9163.n172 a_5396_9163.n6 2.37644
R12918 a_5396_9163.n94 a_5396_9163.n45 2.23844
R12919 a_5396_9163.n246 a_5396_9163.n245 2.2016
R12920 a_5396_9163.n251 a_5396_9163.n250 2.2016
R12921 a_5396_9163.n257 a_5396_9163.n256 2.2016
R12922 a_5396_9163.n263 a_5396_9163.n262 2.2016
R12923 a_5396_9163.n240 a_5396_9163.n239 2.2016
R12924 a_5396_9163.n234 a_5396_9163.n233 2.2016
R12925 a_5396_9163.n228 a_5396_9163.n227 2.2016
R12926 a_5396_9163.n222 a_5396_9163.n221 2.2016
R12927 a_5396_9163.n147 a_5396_9163.n146 2.2016
R12928 a_5396_9163.n152 a_5396_9163.n151 2.2016
R12929 a_5396_9163.n158 a_5396_9163.n157 2.2016
R12930 a_5396_9163.n164 a_5396_9163.n163 2.2016
R12931 a_5396_9163.n179 a_5396_9163.n178 2.2016
R12932 a_5396_9163.n185 a_5396_9163.n184 2.2016
R12933 a_5396_9163.n191 a_5396_9163.n190 2.2016
R12934 a_5396_9163.n197 a_5396_9163.n196 2.2016
R12935 a_5396_9163.n173 a_5396_9163.n172 2.0852
R12936 a_5396_9163.n274 a_5396_9163.n273 1.85726
R12937 a_5396_9163.n281 a_5396_9163.n30 1.83738
R12938 a_5396_9163.n223 a_5396_9163.n138 1.65018
R12939 a_5396_9163.n199 a_5396_9163.n198 1.65018
R12940 a_5396_9163.n96 a_5396_9163.n0 1.65553
R12941 a_5396_9163.n280 a_5396_9163.n3 1.65553
R12942 a_5396_9163.n55 a_5396_9163.n31 1.5005
R12943 a_5396_9163.n203 a_5396_9163.n142 1.5005
R12944 a_5396_9163.n217 a_5396_9163.n216 1.5005
R12945 a_5396_9163.n268 a_5396_9163.n267 1.5005
R12946 a_5396_9163.n174 a_5396_9163.n173 1.5005
R12947 a_5396_9163.n266 a_5396_9163.n265 1.5005
R12948 a_5396_9163.n281 a_5396_9163.n280 1.5005
R12949 a_5396_9163.n102 a_5396_9163.n29 1.5005
R12950 a_5396_9163.n96 a_5396_9163.n95 1.5005
R12951 a_5396_9163.n94 a_5396_9163.n93 1.5005
R12952 a_5396_9163.n283 a_5396_9163.n282 1.5005
R12953 a_5396_9163.n137 a_5396_9163.n136 1.5005
R12954 a_5396_9163.n14 a_5396_9163.t64 1.4705
R12955 a_5396_9163.n14 a_5396_9163.n13 1.4705
R12956 a_5396_9163.n16 a_5396_9163.t43 1.4705
R12957 a_5396_9163.n16 a_5396_9163.n15 1.4705
R12958 a_5396_9163.n24 a_5396_9163.t16 1.4705
R12959 a_5396_9163.n24 a_5396_9163.n23 1.4705
R12960 a_5396_9163.n26 a_5396_9163.t65 1.4705
R12961 a_5396_9163.n26 a_5396_9163.n25 1.4705
R12962 a_5396_9163.n125 a_5396_9163.t53 1.4705
R12963 a_5396_9163.n125 a_5396_9163.n124 1.4705
R12964 a_5396_9163.n127 a_5396_9163.t25 1.4705
R12965 a_5396_9163.n127 a_5396_9163.n126 1.4705
R12966 a_5396_9163.n113 a_5396_9163.t8 1.4705
R12967 a_5396_9163.n113 a_5396_9163.n112 1.4705
R12968 a_5396_9163.n115 a_5396_9163.t15 1.4705
R12969 a_5396_9163.n115 a_5396_9163.n114 1.4705
R12970 a_5396_9163.n42 a_5396_9163.t77 1.4705
R12971 a_5396_9163.n42 a_5396_9163.n41 1.4705
R12972 a_5396_9163.n39 a_5396_9163.t3 1.4705
R12973 a_5396_9163.n39 a_5396_9163.n38 1.4705
R12974 a_5396_9163.n82 a_5396_9163.t26 1.4705
R12975 a_5396_9163.n82 a_5396_9163.n81 1.4705
R12976 a_5396_9163.n84 a_5396_9163.t32 1.4705
R12977 a_5396_9163.n84 a_5396_9163.n83 1.4705
R12978 a_5396_9163.n75 a_5396_9163.t69 1.4705
R12979 a_5396_9163.n75 a_5396_9163.n74 1.4705
R12980 a_5396_9163.n77 a_5396_9163.t74 1.4705
R12981 a_5396_9163.n77 a_5396_9163.n76 1.4705
R12982 a_5396_9163.n63 a_5396_9163.t12 1.4705
R12983 a_5396_9163.n63 a_5396_9163.n62 1.4705
R12984 a_5396_9163.n65 a_5396_9163.t23 1.4705
R12985 a_5396_9163.n65 a_5396_9163.n64 1.4705
R12986 a_5396_9163.n50 a_5396_9163.t62 1.4705
R12987 a_5396_9163.n50 a_5396_9163.n49 1.4705
R12988 a_5396_9163.n52 a_5396_9163.t66 1.4705
R12989 a_5396_9163.n52 a_5396_9163.n51 1.4705
R12990 a_5396_9163.n35 a_5396_9163.t31 1.4705
R12991 a_5396_9163.n35 a_5396_9163.n34 1.4705
R12992 a_5396_9163.n33 a_5396_9163.t45 1.4705
R12993 a_5396_9163.n33 a_5396_9163.n32 1.4705
R12994 a_5396_9163.n99 a_5396_9163.t29 1.4705
R12995 a_5396_9163.n99 a_5396_9163.n98 1.4705
R12996 a_5396_9163.n104 a_5396_9163.t40 1.4705
R12997 a_5396_9163.n104 a_5396_9163.n103 1.4705
R12998 a_5396_9163.n279 a_5396_9163.t36 1.4705
R12999 a_5396_9163.n279 a_5396_9163.n278 1.4705
R13000 a_5396_9163.n277 a_5396_9163.t81 1.4705
R13001 a_5396_9163.n277 a_5396_9163.n276 1.4705
R13002 a_5396_9163.n171 a_5396_9163.t119 1.4705
R13003 a_5396_9163.n171 a_5396_9163.n170 1.4705
R13004 a_5396_9163.n168 a_5396_9163.t130 1.4705
R13005 a_5396_9163.n168 a_5396_9163.n167 1.4705
R13006 a_5396_9163.n243 a_5396_9163.t91 1.4705
R13007 a_5396_9163.n243 a_5396_9163.n242 1.4705
R13008 a_5396_9163.n245 a_5396_9163.t92 1.4705
R13009 a_5396_9163.n245 a_5396_9163.n244 1.4705
R13010 a_5396_9163.n248 a_5396_9163.t121 1.4705
R13011 a_5396_9163.n248 a_5396_9163.n247 1.4705
R13012 a_5396_9163.n250 a_5396_9163.t123 1.4705
R13013 a_5396_9163.n250 a_5396_9163.n249 1.4705
R13014 a_5396_9163.n254 a_5396_9163.t113 1.4705
R13015 a_5396_9163.n254 a_5396_9163.n253 1.4705
R13016 a_5396_9163.n256 a_5396_9163.t114 1.4705
R13017 a_5396_9163.n256 a_5396_9163.n255 1.4705
R13018 a_5396_9163.n260 a_5396_9163.t105 1.4705
R13019 a_5396_9163.n260 a_5396_9163.n259 1.4705
R13020 a_5396_9163.n262 a_5396_9163.t106 1.4705
R13021 a_5396_9163.n262 a_5396_9163.n261 1.4705
R13022 a_5396_9163.n237 a_5396_9163.t124 1.4705
R13023 a_5396_9163.n237 a_5396_9163.n236 1.4705
R13024 a_5396_9163.n239 a_5396_9163.t125 1.4705
R13025 a_5396_9163.n239 a_5396_9163.n238 1.4705
R13026 a_5396_9163.n231 a_5396_9163.t111 1.4705
R13027 a_5396_9163.n231 a_5396_9163.n230 1.4705
R13028 a_5396_9163.n233 a_5396_9163.t112 1.4705
R13029 a_5396_9163.n233 a_5396_9163.n232 1.4705
R13030 a_5396_9163.n225 a_5396_9163.t96 1.4705
R13031 a_5396_9163.n225 a_5396_9163.n224 1.4705
R13032 a_5396_9163.n227 a_5396_9163.t97 1.4705
R13033 a_5396_9163.n227 a_5396_9163.n226 1.4705
R13034 a_5396_9163.n219 a_5396_9163.t126 1.4705
R13035 a_5396_9163.n219 a_5396_9163.n218 1.4705
R13036 a_5396_9163.n221 a_5396_9163.t127 1.4705
R13037 a_5396_9163.n221 a_5396_9163.n220 1.4705
R13038 a_5396_9163.n144 a_5396_9163.t89 1.4705
R13039 a_5396_9163.n144 a_5396_9163.n143 1.4705
R13040 a_5396_9163.n146 a_5396_9163.t88 1.4705
R13041 a_5396_9163.n146 a_5396_9163.n145 1.4705
R13042 a_5396_9163.n149 a_5396_9163.t109 1.4705
R13043 a_5396_9163.n149 a_5396_9163.n148 1.4705
R13044 a_5396_9163.n151 a_5396_9163.t108 1.4705
R13045 a_5396_9163.n151 a_5396_9163.n150 1.4705
R13046 a_5396_9163.n155 a_5396_9163.t99 1.4705
R13047 a_5396_9163.n155 a_5396_9163.n154 1.4705
R13048 a_5396_9163.n157 a_5396_9163.t98 1.4705
R13049 a_5396_9163.n157 a_5396_9163.n156 1.4705
R13050 a_5396_9163.n161 a_5396_9163.t129 1.4705
R13051 a_5396_9163.n161 a_5396_9163.n160 1.4705
R13052 a_5396_9163.n163 a_5396_9163.t128 1.4705
R13053 a_5396_9163.n163 a_5396_9163.n162 1.4705
R13054 a_5396_9163.n176 a_5396_9163.t118 1.4705
R13055 a_5396_9163.n176 a_5396_9163.n175 1.4705
R13056 a_5396_9163.n178 a_5396_9163.t117 1.4705
R13057 a_5396_9163.n178 a_5396_9163.n177 1.4705
R13058 a_5396_9163.n182 a_5396_9163.t104 1.4705
R13059 a_5396_9163.n182 a_5396_9163.n181 1.4705
R13060 a_5396_9163.n184 a_5396_9163.t103 1.4705
R13061 a_5396_9163.n184 a_5396_9163.n183 1.4705
R13062 a_5396_9163.n188 a_5396_9163.t101 1.4705
R13063 a_5396_9163.n188 a_5396_9163.n187 1.4705
R13064 a_5396_9163.n190 a_5396_9163.t100 1.4705
R13065 a_5396_9163.n190 a_5396_9163.n189 1.4705
R13066 a_5396_9163.n194 a_5396_9163.t122 1.4705
R13067 a_5396_9163.n194 a_5396_9163.n193 1.4705
R13068 a_5396_9163.n196 a_5396_9163.t120 1.4705
R13069 a_5396_9163.n196 a_5396_9163.n195 1.4705
R13070 a_5396_9163.n140 a_5396_9163.t95 1.4705
R13071 a_5396_9163.n140 a_5396_9163.n139 1.4705
R13072 a_5396_9163.n271 a_5396_9163.t116 1.4705
R13073 a_5396_9163.n271 a_5396_9163.n270 1.4705
R13074 a_5396_9163.n215 a_5396_9163.t94 1.4705
R13075 a_5396_9163.n215 a_5396_9163.n214 1.4705
R13076 a_5396_9163.n212 a_5396_9163.t115 1.4705
R13077 a_5396_9163.n212 a_5396_9163.n211 1.4705
R13078 a_5396_9163.n201 a_5396_9163.t131 1.4705
R13079 a_5396_9163.n201 a_5396_9163.n200 1.4705
R13080 a_5396_9163.n206 a_5396_9163.t93 1.4705
R13081 a_5396_9163.n206 a_5396_9163.n205 1.4705
R13082 a_5396_9163.n18 a_5396_9163.n17 1.46537
R13083 a_5396_9163.n22 a_5396_9163.n21 1.46537
R13084 a_5396_9163.n28 a_5396_9163.n27 1.46537
R13085 a_5396_9163.n121 a_5396_9163.n120 1.46537
R13086 a_5396_9163.n123 a_5396_9163.n122 1.46537
R13087 a_5396_9163.n129 a_5396_9163.n128 1.46537
R13088 a_5396_9163.n133 a_5396_9163.n132 1.46537
R13089 a_5396_9163.n117 a_5396_9163.n116 1.46537
R13090 a_5396_9163.n86 a_5396_9163.n85 1.46537
R13091 a_5396_9163.n90 a_5396_9163.n89 1.46537
R13092 a_5396_9163.n79 a_5396_9163.n78 1.46537
R13093 a_5396_9163.n73 a_5396_9163.n72 1.46537
R13094 a_5396_9163.n69 a_5396_9163.n68 1.46537
R13095 a_5396_9163.n67 a_5396_9163.n66 1.46537
R13096 a_5396_9163.n61 a_5396_9163.n60 1.46537
R13097 a_5396_9163.n54 a_5396_9163.n53 1.46537
R13098 a_5396_9163.n252 a_5396_9163.n251 1.46537
R13099 a_5396_9163.n258 a_5396_9163.n257 1.46537
R13100 a_5396_9163.n264 a_5396_9163.n263 1.46537
R13101 a_5396_9163.n241 a_5396_9163.n240 1.46537
R13102 a_5396_9163.n235 a_5396_9163.n234 1.46537
R13103 a_5396_9163.n229 a_5396_9163.n228 1.46537
R13104 a_5396_9163.n223 a_5396_9163.n222 1.46537
R13105 a_5396_9163.n153 a_5396_9163.n152 1.46537
R13106 a_5396_9163.n159 a_5396_9163.n158 1.46537
R13107 a_5396_9163.n165 a_5396_9163.n164 1.46537
R13108 a_5396_9163.n180 a_5396_9163.n179 1.46537
R13109 a_5396_9163.n186 a_5396_9163.n185 1.46537
R13110 a_5396_9163.n192 a_5396_9163.n191 1.46537
R13111 a_5396_9163.n198 a_5396_9163.n197 1.46537
R13112 a_5396_9163.n285 a_5396_9163.n284 1.46535
R13113 a_5396_9163.n135 a_5396_9163.n134 1.46535
R13114 a_5396_9163.n92 a_5396_9163.n91 1.46535
R13115 a_5396_9163.n57 a_5396_9163.n56 1.46535
R13116 a_5396_9163.n40 a_5396_9163.n37 1.27228
R13117 a_5396_9163.n67 a_5396_9163.n61 1.27228
R13118 a_5396_9163.n69 a_5396_9163.n67 1.27228
R13119 a_5396_9163.n79 a_5396_9163.n73 1.27228
R13120 a_5396_9163.n90 a_5396_9163.n86 1.27228
R13121 a_5396_9163.n107 a_5396_9163.n105 1.27228
R13122 a_5396_9163.n133 a_5396_9163.n129 1.27228
R13123 a_5396_9163.n129 a_5396_9163.n123 1.27228
R13124 a_5396_9163.n121 a_5396_9163.n28 1.27228
R13125 a_5396_9163.n22 a_5396_9163.n18 1.27228
R13126 a_5396_9163.n229 a_5396_9163.n223 1.27228
R13127 a_5396_9163.n241 a_5396_9163.n235 1.27228
R13128 a_5396_9163.n264 a_5396_9163.n258 1.27228
R13129 a_5396_9163.n198 a_5396_9163.n192 1.27228
R13130 a_5396_9163.n186 a_5396_9163.n180 1.27228
R13131 a_5396_9163.n165 a_5396_9163.n159 1.27228
R13132 a_5396_9163.n272 a_5396_9163.n269 1.27228
R13133 a_5396_9163.n207 a_5396_9163.n204 1.27228
R13134 a_5396_9163.n267 a_5396_9163.n30 1.25341
R13135 a_5396_9163.n275 a_5396_9163.n274 1.23151
R13136 a_5396_9163.n45 a_5396_9163.n44 1.01873
R13137 a_5396_9163.n102 a_5396_9163.n101 1.01873
R13138 a_5396_9163.n97 a_5396_9163.n31 0.778574
R13139 a_5396_9163.n275 a_5396_9163.n137 0.778574
R13140 a_5396_9163.n95 a_5396_9163.n94 0.778574
R13141 a_5396_9163.n282 a_5396_9163.n281 0.778574
R13142 a_5396_9163.n137 a_5396_9163.n108 0.738439
R13143 a_5396_9163.n282 a_5396_9163.n29 0.738439
R13144 a_5396_9163.n273 a_5396_9163.n138 0.737223
R13145 a_5396_9163.n208 a_5396_9163.n199 0.737223
R13146 a_5396_9163.n267 a_5396_9163.n266 0.737223
R13147 a_5396_9163.n173 a_5396_9163.n142 0.737223
R13148 a_5396_9163.n209 a_5396_9163.n208 0.725061
R13149 a_5396_9163.n217 a_5396_9163.n142 0.725061
R13150 a_5396_9163.n57 a_5396_9163.n55 0.699581
R13151 a_5396_9163.n93 a_5396_9163.n92 0.699581
R13152 a_5396_9163.n136 a_5396_9163.n135 0.699581
R13153 a_5396_9163.n284 a_5396_9163.n283 0.699581
R13154 a_5396_9163.n209 a_5396_9163.n138 0.585196
R13155 a_5396_9163.n266 a_5396_9163.n217 0.585196
R13156 a_5396_9163.n55 a_5396_9163.n54 0.557791
R13157 a_5396_9163.n93 a_5396_9163.n79 0.557791
R13158 a_5396_9163.n136 a_5396_9163.n117 0.557791
R13159 a_5396_9163.n283 a_5396_9163.n28 0.557791
R13160 a_5396_9163.n108 a_5396_9163.n97 0.530466
R13161 a_5396_9163.n95 a_5396_9163.n29 0.530466
R13162 a_5396_9163.n265 a_5396_9163.n264 0.150184
R13163 a_5396_9163.n174 a_5396_9163.n165 0.150184
R13164 a_5396_9163.n1 a_5396_9163.n2 1.27228
R13165 a_5396_9163.n96 a_5396_9163.n1 7.30549
R13166 a_5396_9163.t71 a_5396_9163.n0 6.96214
R13167 a_5396_9163.n4 a_5396_9163.n5 1.27228
R13168 a_5396_9163.n280 a_5396_9163.n4 7.30549
R13169 a_5396_9163.t58 a_5396_9163.n3 6.96214
R13170 a_5396_9163.n10 a_5396_9163.n11 1.26457
R13171 a_5396_9163.n216 a_5396_9163.n10 6.59229
R13172 a_5396_9163.n215 a_5396_9163.n9 5.10549
R13173 a_5396_9163.n7 a_5396_9163.n8 1.26457
R13174 a_5396_9163.n172 a_5396_9163.n7 6.59229
R13175 a_5396_9163.n171 a_5396_9163.n6 5.10549
R13176 VOUT.n35 VOUT.n23 7.94229
R13177 VOUT.n104 VOUT.n101 7.94229
R13178 VOUT.n98 VOUT.n90 7.169
R13179 VOUT.n191 VOUT.n190 7.169
R13180 VOUT.n162 VOUT.t16 6.96668
R13181 VOUT.n10 VOUT.t67 6.82564
R13182 VOUT.n95 VOUT.t89 6.82564
R13183 VOUT.n186 VOUT.n185 5.85326
R13184 VOUT.n186 VOUT.n184 5.84661
R13185 VOUT.n22 VOUT.n21 5.69423
R13186 VOUT.n37 VOUT.n36 5.69423
R13187 VOUT.n18 VOUT.n17 5.69423
R13188 VOUT.n106 VOUT.n105 5.69423
R13189 VOUT.n22 VOUT.n20 5.49558
R13190 VOUT.n18 VOUT.n16 5.49558
R13191 VOUT.n12 VOUT.n11 4.61332
R13192 VOUT.n193 VOUT.n192 4.61332
R13193 VOUT.n97 VOUT.n96 4.61332
R13194 VOUT.n89 VOUT.n87 4.61332
R13195 VOUT.n85 VOUT.n81 4.61332
R13196 VOUT.n164 VOUT.n163 4.61332
R13197 VOUT.n3 VOUT.n2 4.61332
R13198 VOUT.n11 VOUT.n10 4.60571
R13199 VOUT.n192 VOUT.n191 4.60571
R13200 VOUT.n96 VOUT.n95 4.60571
R13201 VOUT.n90 VOUT.n89 4.60571
R13202 VOUT.n86 VOUT.n85 4.60571
R13203 VOUT.n163 VOUT.n162 4.60571
R13204 VOUT.n194 VOUT.n2 4.60571
R13205 VOUT.n84 VOUT.n80 4.5005
R13206 VOUT.n88 VOUT.n79 4.5005
R13207 VOUT.n94 VOUT.n91 4.5005
R13208 VOUT.n161 VOUT.n158 4.5005
R13209 VOUT.n5 VOUT.n4 4.5005
R13210 VOUT.n9 VOUT.n6 4.5005
R13211 VOUT.n196 VOUT.n195 4.5005
R13212 VOUT.n5 VOUT.t82 4.22462
R13213 VOUT.n88 VOUT.t48 4.22462
R13214 VOUT.n35 VOUT.n34 4.22423
R13215 VOUT.n104 VOUT.n103 4.22423
R13216 VOUT.n177 VOUT.n176 4.21195
R13217 VOUT.n179 VOUT.t6 4.21195
R13218 VOUT.n64 VOUT.t73 4.05054
R13219 VOUT.n73 VOUT.n72 4.05054
R13220 VOUT.n75 VOUT.t75 4.05054
R13221 VOUT.n56 VOUT.n55 4.05054
R13222 VOUT.n52 VOUT.t34 4.05054
R13223 VOUT.n44 VOUT.n43 4.05054
R13224 VOUT.n40 VOUT.t40 4.05054
R13225 VOUT.n26 VOUT.n25 4.05054
R13226 VOUT.n117 VOUT.t47 4.05054
R13227 VOUT.n126 VOUT.n125 4.05054
R13228 VOUT.n128 VOUT.t22 4.05054
R13229 VOUT.n139 VOUT.n138 4.05054
R13230 VOUT.n141 VOUT.t60 4.05054
R13231 VOUT.n151 VOUT.n150 4.05054
R13232 VOUT.n153 VOUT.t33 4.05054
R13233 VOUT.n110 VOUT.n109 4.05054
R13234 VOUT.n177 VOUT.n175 4.03668
R13235 VOUT.n179 VOUT.t13 4.03668
R13236 VOUT.n64 VOUT.t69 3.87765
R13237 VOUT.n73 VOUT.n71 3.87765
R13238 VOUT.n75 VOUT.t72 3.87765
R13239 VOUT.n56 VOUT.n54 3.87765
R13240 VOUT.n52 VOUT.t32 3.87765
R13241 VOUT.n44 VOUT.n42 3.87765
R13242 VOUT.n40 VOUT.t39 3.87765
R13243 VOUT.n26 VOUT.n24 3.87765
R13244 VOUT.n117 VOUT.t49 3.87765
R13245 VOUT.n126 VOUT.n124 3.87765
R13246 VOUT.n128 VOUT.t23 3.87765
R13247 VOUT.n139 VOUT.n137 3.87765
R13248 VOUT.n141 VOUT.t61 3.87765
R13249 VOUT.n151 VOUT.n149 3.87765
R13250 VOUT.n153 VOUT.t35 3.87765
R13251 VOUT.n110 VOUT.n108 3.87765
R13252 VOUT.n182 VOUT.n164 3.81532
R13253 VOUT.n189 VOUT.n188 3.544
R13254 VOUT.n188 VOUT.n157 3.48165
R13255 VOUT.n38 VOUT.n37 3.25667
R13256 VOUT.n161 VOUT.n160 3.12366
R13257 VOUT.n81 VOUT.n14 3.01925
R13258 VOUT.n157 VOUT.n3 3.01925
R13259 VOUT.n174 VOUT.n173 2.95195
R13260 VOUT.n169 VOUT.n168 2.95195
R13261 VOUT.n174 VOUT.n171 2.77668
R13262 VOUT.n169 VOUT.n166 2.77668
R13263 VOUT.n9 VOUT.n8 2.75462
R13264 VOUT.n94 VOUT.n93 2.75462
R13265 VOUT.n84 VOUT.n83 2.75462
R13266 VOUT.n32 VOUT.n26 2.73714
R13267 VOUT.n116 VOUT.n110 2.73714
R13268 VOUT.n70 VOUT.n64 2.73672
R13269 VOUT.n123 VOUT.n117 2.73672
R13270 VOUT.n178 VOUT.n174 2.71872
R13271 VOUT.n57 VOUT.n53 2.60203
R13272 VOUT.n142 VOUT.n140 2.60203
R13273 VOUT.n69 VOUT.n68 2.58054
R13274 VOUT.n62 VOUT.n61 2.58054
R13275 VOUT.n50 VOUT.n49 2.58054
R13276 VOUT.n31 VOUT.n30 2.58054
R13277 VOUT.n122 VOUT.n121 2.58054
R13278 VOUT.n135 VOUT.n134 2.58054
R13279 VOUT.n147 VOUT.n146 2.58054
R13280 VOUT.n115 VOUT.n114 2.58054
R13281 VOUT.n180 VOUT.n178 2.56118
R13282 VOUT.n187 VOUT.n186 2.54573
R13283 VOUT.n45 VOUT.n41 2.53418
R13284 VOUT.n76 VOUT.n74 2.53418
R13285 VOUT.n154 VOUT.n152 2.53418
R13286 VOUT.n129 VOUT.n127 2.53418
R13287 VOUT.n107 VOUT.n106 2.51873
R13288 VOUT.n69 VOUT.n66 2.40765
R13289 VOUT.n62 VOUT.n59 2.40765
R13290 VOUT.n50 VOUT.n47 2.40765
R13291 VOUT.n31 VOUT.n28 2.40765
R13292 VOUT.n122 VOUT.n119 2.40765
R13293 VOUT.n135 VOUT.n132 2.40765
R13294 VOUT.n147 VOUT.n144 2.40765
R13295 VOUT.n115 VOUT.n112 2.40765
R13296 VOUT.n78 VOUT.n23 2.23844
R13297 VOUT VOUT.n1 2.05949
R13298 VOUT.n181 VOUT.n169 2.00466
R13299 VOUT.n98 VOUT.n97 1.51925
R13300 VOUT.n190 VOUT.n12 1.51925
R13301 VOUT.n156 VOUT.n155 1.5005
R13302 VOUT.n39 VOUT.n38 1.5005
R13303 VOUT.n182 VOUT.n181 1.5005
R13304 VOUT.n130 VOUT.n13 1.5005
R13305 VOUT.n101 VOUT.n100 1.5005
R13306 VOUT.n99 VOUT.n98 1.5005
R13307 VOUT.n78 VOUT.n77 1.5005
R13308 VOUT.n190 VOUT.n189 1.5005
R13309 VOUT.n1 VOUT.t43 1.4705
R13310 VOUT.n1 VOUT.n0 1.4705
R13311 VOUT.n8 VOUT.t30 1.4705
R13312 VOUT.n8 VOUT.n7 1.4705
R13313 VOUT.n20 VOUT.t63 1.4705
R13314 VOUT.n20 VOUT.n19 1.4705
R13315 VOUT.n34 VOUT.t21 1.4705
R13316 VOUT.n34 VOUT.n33 1.4705
R13317 VOUT.n66 VOUT.t29 1.4705
R13318 VOUT.n66 VOUT.n65 1.4705
R13319 VOUT.n68 VOUT.t31 1.4705
R13320 VOUT.n68 VOUT.n67 1.4705
R13321 VOUT.n59 VOUT.t53 1.4705
R13322 VOUT.n59 VOUT.n58 1.4705
R13323 VOUT.n61 VOUT.t54 1.4705
R13324 VOUT.n61 VOUT.n60 1.4705
R13325 VOUT.n47 VOUT.t100 1.4705
R13326 VOUT.n47 VOUT.n46 1.4705
R13327 VOUT.n49 VOUT.t102 1.4705
R13328 VOUT.n49 VOUT.n48 1.4705
R13329 VOUT.n28 VOUT.t92 1.4705
R13330 VOUT.n28 VOUT.n27 1.4705
R13331 VOUT.n30 VOUT.t94 1.4705
R13332 VOUT.n30 VOUT.n29 1.4705
R13333 VOUT.n93 VOUT.t95 1.4705
R13334 VOUT.n93 VOUT.n92 1.4705
R13335 VOUT.n83 VOUT.t50 1.4705
R13336 VOUT.n83 VOUT.n82 1.4705
R13337 VOUT.n16 VOUT.t76 1.4705
R13338 VOUT.n16 VOUT.n15 1.4705
R13339 VOUT.n103 VOUT.t84 1.4705
R13340 VOUT.n103 VOUT.n102 1.4705
R13341 VOUT.n119 VOUT.t37 1.4705
R13342 VOUT.n119 VOUT.n118 1.4705
R13343 VOUT.n121 VOUT.t36 1.4705
R13344 VOUT.n121 VOUT.n120 1.4705
R13345 VOUT.n132 VOUT.t81 1.4705
R13346 VOUT.n132 VOUT.n131 1.4705
R13347 VOUT.n134 VOUT.t79 1.4705
R13348 VOUT.n134 VOUT.n133 1.4705
R13349 VOUT.n144 VOUT.t27 1.4705
R13350 VOUT.n144 VOUT.n143 1.4705
R13351 VOUT.n146 VOUT.t26 1.4705
R13352 VOUT.n146 VOUT.n145 1.4705
R13353 VOUT.n112 VOUT.t70 1.4705
R13354 VOUT.n112 VOUT.n111 1.4705
R13355 VOUT.n114 VOUT.t68 1.4705
R13356 VOUT.n114 VOUT.n113 1.4705
R13357 VOUT.n70 VOUT.n69 1.46537
R13358 VOUT.n74 VOUT.n73 1.46537
R13359 VOUT.n63 VOUT.n62 1.46537
R13360 VOUT.n57 VOUT.n56 1.46537
R13361 VOUT.n53 VOUT.n52 1.46537
R13362 VOUT.n51 VOUT.n50 1.46537
R13363 VOUT.n45 VOUT.n44 1.46537
R13364 VOUT.n32 VOUT.n31 1.46537
R13365 VOUT.n123 VOUT.n122 1.46537
R13366 VOUT.n127 VOUT.n126 1.46537
R13367 VOUT.n136 VOUT.n135 1.46537
R13368 VOUT.n140 VOUT.n139 1.46537
R13369 VOUT.n142 VOUT.n141 1.46537
R13370 VOUT.n148 VOUT.n147 1.46537
R13371 VOUT.n152 VOUT.n151 1.46537
R13372 VOUT.n116 VOUT.n115 1.46537
R13373 VOUT.n178 VOUT.n177 1.46537
R13374 VOUT.n76 VOUT.n75 1.46535
R13375 VOUT.n41 VOUT.n40 1.46535
R13376 VOUT.n129 VOUT.n128 1.46535
R13377 VOUT.n154 VOUT.n153 1.46535
R13378 VOUT.n180 VOUT.n179 1.46535
R13379 VOUT.n37 VOUT.n35 1.27228
R13380 VOUT.n51 VOUT.n45 1.27228
R13381 VOUT.n53 VOUT.n51 1.27228
R13382 VOUT.n63 VOUT.n57 1.27228
R13383 VOUT.n74 VOUT.n70 1.27228
R13384 VOUT.n106 VOUT.n104 1.27228
R13385 VOUT.n152 VOUT.n148 1.27228
R13386 VOUT.n148 VOUT.n142 1.27228
R13387 VOUT.n140 VOUT.n136 1.27228
R13388 VOUT.n127 VOUT.n123 1.27228
R13389 VOUT.n184 VOUT.t11 1.2605
R13390 VOUT.n184 VOUT.n183 1.2605
R13391 VOUT.n171 VOUT.t15 1.2605
R13392 VOUT.n171 VOUT.n170 1.2605
R13393 VOUT.n173 VOUT.t8 1.2605
R13394 VOUT.n173 VOUT.n172 1.2605
R13395 VOUT.n166 VOUT.t14 1.2605
R13396 VOUT.n166 VOUT.n165 1.2605
R13397 VOUT.n168 VOUT.t7 1.2605
R13398 VOUT.n168 VOUT.n167 1.2605
R13399 VOUT.n160 VOUT.t17 1.2605
R13400 VOUT.n160 VOUT.n159 1.2605
R13401 VOUT.n188 VOUT.n187 1.25797
R13402 VOUT.n23 VOUT.n22 1.01873
R13403 VOUT.n101 VOUT.n18 1.01873
R13404 VOUT.n87 VOUT.n86 0.9995
R13405 VOUT.n194 VOUT.n193 0.9995
R13406 VOUT.n38 VOUT.n14 0.778574
R13407 VOUT.n157 VOUT.n156 0.778574
R13408 VOUT.n99 VOUT.n78 0.778574
R13409 VOUT.n189 VOUT.n13 0.778574
R13410 VOUT.n156 VOUT.n107 0.738439
R13411 VOUT.n187 VOUT.n182 0.738439
R13412 VOUT.n100 VOUT.n13 0.738439
R13413 VOUT.n41 VOUT.n39 0.699581
R13414 VOUT.n77 VOUT.n76 0.699581
R13415 VOUT.n155 VOUT.n154 0.699581
R13416 VOUT.n130 VOUT.n129 0.699581
R13417 VOUT.n181 VOUT.n180 0.699581
R13418 VOUT VOUT.n196 0.695632
R13419 VOUT.n39 VOUT.n32 0.557791
R13420 VOUT.n77 VOUT.n63 0.557791
R13421 VOUT.n155 VOUT.n116 0.557791
R13422 VOUT.n136 VOUT.n130 0.557791
R13423 VOUT.n107 VOUT.n14 0.530466
R13424 VOUT.n100 VOUT.n99 0.530466
R13425 VOUT.n81 VOUT.n80 0.14
R13426 VOUT.n86 VOUT.n80 0.14
R13427 VOUT.n87 VOUT.n79 0.14
R13428 VOUT.n90 VOUT.n79 0.14
R13429 VOUT.n97 VOUT.n91 0.14
R13430 VOUT.n95 VOUT.n91 0.14
R13431 VOUT.n164 VOUT.n158 0.14
R13432 VOUT.n162 VOUT.n158 0.14
R13433 VOUT.n195 VOUT.n3 0.14
R13434 VOUT.n195 VOUT.n194 0.14
R13435 VOUT.n193 VOUT.n4 0.14
R13436 VOUT.n191 VOUT.n4 0.14
R13437 VOUT.n12 VOUT.n6 0.14
R13438 VOUT.n10 VOUT.n6 0.14
R13439 VOUT.n11 VOUT.n9 0.00168421
R13440 VOUT.n192 VOUT.n5 0.00168421
R13441 VOUT.n96 VOUT.n94 0.00168421
R13442 VOUT.n89 VOUT.n88 0.00168421
R13443 VOUT.n85 VOUT.n84 0.00168421
R13444 VOUT.n163 VOUT.n161 0.00168421
R13445 VOUT.n196 VOUT.n2 0.00168421
R13446 a_n11737_n14973.n337 a_n11737_n14973.t4 10.621
R13447 a_n11737_n14973.n333 a_n11737_n14973.t35 10.621
R13448 a_n11737_n14973.n344 a_n11737_n14973.n330 10.3121
R13449 a_n11737_n14973.n339 a_n11737_n14973.t79 10.3044
R13450 a_n11737_n14973.n335 a_n11737_n14973.t6 10.3044
R13451 a_n11737_n14973.n338 a_n11737_n14973.t97 9.9994
R13452 a_n11737_n14973.n334 a_n11737_n14973.t2 9.9994
R13453 a_n11737_n14973.n337 a_n11737_n14973.t0 9.999
R13454 a_n11737_n14973.n333 a_n11737_n14973.t48 9.999
R13455 a_n11737_n14973.n228 a_n11737_n14973.t54 8.33806
R13456 a_n11737_n14973.n323 a_n11737_n14973.t95 8.3366
R13457 a_n11737_n14973.n282 a_n11737_n14973.t78 8.26493
R13458 a_n11737_n14973.n96 a_n11737_n14973.t71 8.35715
R13459 a_n11737_n14973.n43 a_n11737_n14973.t101 8.06917
R13460 a_n11737_n14973.n55 a_n11737_n14973.t69 8.06917
R13461 a_n11737_n14973.n122 a_n11737_n14973.t92 8.06917
R13462 a_n11737_n14973.n31 a_n11737_n14973.t77 8.06917
R13463 a_n11737_n14973.n132 a_n11737_n14973.t106 8.06917
R13464 a_n11737_n14973.n50 a_n11737_n14973.t55 8.06917
R13465 a_n11737_n14973.n57 a_n11737_n14973.t31 8.06917
R13466 a_n11737_n14973.n17 a_n11737_n14973.t44 8.06917
R13467 a_n11737_n14973.n78 a_n11737_n14973.t33 8.06917
R13468 a_n11737_n14973.n28 a_n11737_n14973.t86 8.06917
R13469 a_n11737_n14973.n133 a_n11737_n14973.t32 8.06917
R13470 a_n11737_n14973.n9 a_n11737_n14973.t47 8.06917
R13471 a_n11737_n14973.n8 a_n11737_n14973.t34 8.06917
R13472 a_n11737_n14973.n174 a_n11737_n14973.t45 8.06917
R13473 a_n11737_n14973.n6 a_n11737_n14973.t81 8.06917
R13474 a_n11737_n14973.n5 a_n11737_n14973.t57 8.06917
R13475 a_n11737_n14973.n179 a_n11737_n14973.t80 8.06917
R13476 a_n11737_n14973.n40 a_n11737_n14973.t68 8.06917
R13477 a_n11737_n14973.n93 a_n11737_n14973.t76 8.06917
R13478 a_n11737_n14973.n75 a_n11737_n14973.t49 8.06917
R13479 a_n11737_n14973.n61 a_n11737_n14973.t75 8.06917
R13480 a_n11737_n14973.n34 a_n11737_n14973.t30 8.06917
R13481 a_n11737_n14973.n90 a_n11737_n14973.t82 8.06917
R13482 a_n11737_n14973.n2 a_n11737_n14973.t102 8.06917
R13483 a_n11737_n14973.n86 a_n11737_n14973.t84 8.06917
R13484 a_n11737_n14973.n71 a_n11737_n14973.t53 8.06917
R13485 a_n11737_n14973.n65 a_n11737_n14973.t83 8.06917
R13486 a_n11737_n14973.n125 a_n11737_n14973.t66 8.06917
R13487 a_n11737_n14973.n23 a_n11737_n14973.t50 8.06917
R13488 a_n11737_n14973.n167 a_n11737_n14973.t65 8.06917
R13489 a_n11737_n14973.n128 a_n11737_n14973.t104 8.06917
R13490 a_n11737_n14973.n20 a_n11737_n14973.t88 8.06917
R13491 a_n11737_n14973.n156 a_n11737_n14973.t103 8.06917
R13492 a_n11737_n14973.n82 a_n11737_n14973.t41 8.06917
R13493 a_n11737_n14973.n68 a_n11737_n14973.t58 8.06917
R13494 a_n11737_n14973.n108 a_n11737_n14973.t105 8.06917
R13495 a_n11737_n14973.n97 a_n11737_n14973.t72 8.06917
R13496 a_n11737_n14973.n263 a_n11737_n14973.t93 8.06917
R13497 a_n11737_n14973.n252 a_n11737_n14973.t85 8.06917
R13498 a_n11737_n14973.n251 a_n11737_n14973.t60 8.06917
R13499 a_n11737_n14973.n250 a_n11737_n14973.t87 8.06917
R13500 a_n11737_n14973.n95 a_n11737_n14973.t42 8.06917
R13501 a_n11737_n14973.n243 a_n11737_n14973.t70 8.06917
R13502 a_n11737_n14973.n112 a_n11737_n14973.t61 8.06917
R13503 a_n11737_n14973.n229 a_n11737_n14973.t40 8.06917
R13504 a_n11737_n14973.n235 a_n11737_n14973.t36 8.06917
R13505 a_n11737_n14973.n236 a_n11737_n14973.t96 8.06917
R13506 a_n11737_n14973.n237 a_n11737_n14973.t37 8.06917
R13507 a_n11737_n14973.n109 a_n11737_n14973.t74 8.06917
R13508 a_n11737_n14973.n100 a_n11737_n14973.t46 8.06917
R13509 a_n11737_n14973.n271 a_n11737_n14973.t73 8.06917
R13510 a_n11737_n14973.n322 a_n11737_n14973.t63 8.06917
R13511 a_n11737_n14973.n118 a_n11737_n14973.t94 8.06917
R13512 a_n11737_n14973.n320 a_n11737_n14973.t52 8.06917
R13513 a_n11737_n14973.n319 a_n11737_n14973.t38 8.06917
R13514 a_n11737_n14973.n318 a_n11737_n14973.t51 8.06917
R13515 a_n11737_n14973.n316 a_n11737_n14973.t43 8.06917
R13516 a_n11737_n14973.n309 a_n11737_n14973.t98 8.06917
R13517 a_n11737_n14973.n115 a_n11737_n14973.t39 8.06917
R13518 a_n11737_n14973.n304 a_n11737_n14973.t100 8.06917
R13519 a_n11737_n14973.n101 a_n11737_n14973.t67 8.06917
R13520 a_n11737_n14973.n119 a_n11737_n14973.t99 8.06917
R13521 a_n11737_n14973.n293 a_n11737_n14973.t90 8.06917
R13522 a_n11737_n14973.n292 a_n11737_n14973.t64 8.06917
R13523 a_n11737_n14973.n291 a_n11737_n14973.t89 8.06917
R13524 a_n11737_n14973.n278 a_n11737_n14973.t91 8.06917
R13525 a_n11737_n14973.n281 a_n11737_n14973.t56 8.06917
R13526 a_n11737_n14973.t29 a_n11737_n14973.n372 6.49245
R13527 a_n11737_n14973.n145 a_n11737_n14973.n142 6.49245
R13528 a_n11737_n14973.n140 a_n11737_n14973.n352 6.50349
R13529 a_n11737_n14973.n342 a_n11737_n14973.n341 5.70664
R13530 a_n11737_n14973.n332 a_n11737_n14973.t7 5.23357
R13531 a_n11737_n14973.n146 a_n11737_n14973.t18 5.22068
R13532 a_n11737_n14973.n332 a_n11737_n14973.n331 5.15078
R13533 a_n11737_n14973.n342 a_n11737_n14973.t1 4.6582
R13534 a_n11737_n14973.n84 a_n11737_n14973.n69 2.0194
R13535 a_n11737_n14973.n182 a_n11737_n14973.n123 2.42484
R13536 a_n11737_n14973.n123 a_n11737_n14973.n181 2.4256
R13537 a_n11737_n14973.n110 a_n11737_n14973.n109 2.25048
R13538 a_n11737_n14973.n115 a_n11737_n14973.n113 2.25048
R13539 a_n11737_n14973.n136 a_n11737_n14973.n348 3.76239
R13540 a_n11737_n14973.n137 a_n11737_n14973.n346 5.23239
R13541 a_n11737_n14973.n359 a_n11737_n14973.n358 4.60825
R13542 a_n11737_n14973.n354 a_n11737_n14973.n140 3.76239
R13543 a_n11737_n14973.n10 a_n11737_n14973.n9 1.44552
R13544 a_n11737_n14973.n7 a_n11737_n14973.n6 1.44552
R13545 a_n11737_n14973.n126 a_n11737_n14973.n125 2.22591
R13546 a_n11737_n14973.n129 a_n11737_n14973.n128 2.22591
R13547 a_n11737_n14973.n85 a_n11737_n14973.n163 4.51491
R13548 a_n11737_n14973.n220 a_n11737_n14973.n219 4.51075
R13549 a_n11737_n14973.n62 a_n11737_n14973.n61 2.21906
R13550 a_n11737_n14973.n66 a_n11737_n14973.n65 2.21906
R13551 a_n11737_n14973.n34 a_n11737_n14973.n35 2.21826
R13552 a_n11737_n14973.n40 a_n11737_n14973.n39 2.21826
R13553 a_n11737_n14973.n358 a_n11737_n14973.n345 4.50168
R13554 a_n11737_n14973.n356 a_n11737_n14973.n355 4.5005
R13555 a_n11737_n14973.n139 a_n11737_n14973.n138 2.24327
R13556 a_n11737_n14973.n12 a_n11737_n14973.n5 2.21666
R13557 a_n11737_n14973.n11 a_n11737_n14973.n178 4.5005
R13558 a_n11737_n14973.n188 a_n11737_n14973.n187 4.5005
R13559 a_n11737_n14973.n14 a_n11737_n14973.n8 2.21666
R13560 a_n11737_n14973.n13 a_n11737_n14973.n173 4.5005
R13561 a_n11737_n14973.n206 a_n11737_n14973.n205 4.5005
R13562 a_n11737_n14973.n198 a_n11737_n14973.n197 4.5005
R13563 a_n11737_n14973.n78 a_n11737_n14973.n79 2.21666
R13564 a_n11737_n14973.n195 a_n11737_n14973.n27 4.5005
R13565 a_n11737_n14973.n28 a_n11737_n14973.n25 2.21666
R13566 a_n11737_n14973.n26 a_n11737_n14973.n194 4.5005
R13567 a_n11737_n14973.n193 a_n11737_n14973.n133 4.5005
R13568 a_n11737_n14973.n192 a_n11737_n14973.n191 4.5005
R13569 a_n11737_n14973.n51 a_n11737_n14973.n50 2.21666
R13570 a_n11737_n14973.n200 a_n11737_n14973.n49 4.5005
R13571 a_n11737_n14973.n202 a_n11737_n14973.n201 4.5005
R13572 a_n11737_n14973.n58 a_n11737_n14973.n57 2.21666
R13573 a_n11737_n14973.n16 a_n11737_n14973.n175 4.5005
R13574 a_n11737_n14973.n18 a_n11737_n14973.n17 2.21666
R13575 a_n11737_n14973.n0 a_n11737_n14973.n1 0.0657695
R13576 a_n11737_n14973.n30 a_n11737_n14973.n210 4.5005
R13577 a_n11737_n14973.n32 a_n11737_n14973.n31 2.21666
R13578 a_n11737_n14973.n131 a_n11737_n14973.n209 4.5005
R13579 a_n11737_n14973.n132 a_n11737_n14973.n208 4.5005
R13580 a_n11737_n14973.n212 a_n11737_n14973.n207 4.5005
R13581 a_n11737_n14973.n44 a_n11737_n14973.n43 2.21666
R13582 a_n11737_n14973.n42 a_n11737_n14973.n185 4.5005
R13583 a_n11737_n14973.n184 a_n11737_n14973.n54 4.5005
R13584 a_n11737_n14973.n55 a_n11737_n14973.n52 2.21666
R13585 a_n11737_n14973.n53 a_n11737_n14973.n182 4.5005
R13586 a_n11737_n14973.n123 a_n11737_n14973.n122 0.0107891
R13587 a_n11737_n14973.n127 a_n11737_n14973.n162 4.5005
R13588 a_n11737_n14973.n21 a_n11737_n14973.n20 2.21666
R13589 a_n11737_n14973.n19 a_n11737_n14973.n155 4.5005
R13590 a_n11737_n14973.n161 a_n11737_n14973.n160 4.5005
R13591 a_n11737_n14973.n124 a_n11737_n14973.n170 4.5005
R13592 a_n11737_n14973.n24 a_n11737_n14973.n23 2.21666
R13593 a_n11737_n14973.n22 a_n11737_n14973.n166 4.5005
R13594 a_n11737_n14973.n169 a_n11737_n14973.n168 4.5005
R13595 a_n11737_n14973.n65 a_n11737_n14973.n67 2.21666
R13596 a_n11737_n14973.n64 a_n11737_n14973.n107 4.5005
R13597 a_n11737_n14973.n71 a_n11737_n14973.n73 2.21666
R13598 a_n11737_n14973.n70 a_n11737_n14973.n105 4.5005
R13599 a_n11737_n14973.n86 a_n11737_n14973.n88 2.21666
R13600 a_n11737_n14973.n219 a_n11737_n14973.n218 4.5005
R13601 a_n11737_n14973.n2 a_n11737_n14973.n3 2.21666
R13602 a_n11737_n14973.n90 a_n11737_n14973.n92 2.21666
R13603 a_n11737_n14973.n89 a_n11737_n14973.n102 4.5005
R13604 a_n11737_n14973.n164 a_n11737_n14973.n120 4.5005
R13605 a_n11737_n14973.n36 a_n11737_n14973.n34 2.21666
R13606 a_n11737_n14973.n61 a_n11737_n14973.n63 2.21666
R13607 a_n11737_n14973.n60 a_n11737_n14973.n106 4.5005
R13608 a_n11737_n14973.n75 a_n11737_n14973.n77 2.21666
R13609 a_n11737_n14973.n74 a_n11737_n14973.n104 4.5005
R13610 a_n11737_n14973.n68 a_n11737_n14973.n69 0.0231698
R13611 a_n11737_n14973.n82 a_n11737_n14973.n84 2.21666
R13612 a_n11737_n14973.n157 a_n11737_n14973.n81 4.5005
R13613 a_n11737_n14973.n121 a_n11737_n14973.n158 4.5005
R13614 a_n11737_n14973.n41 a_n11737_n14973.n40 2.21666
R13615 a_n11737_n14973.n83 a_n11737_n14973.n82 2.21666
R13616 a_n11737_n14973.n81 a_n11737_n14973.n103 4.5005
R13617 a_n11737_n14973.n38 a_n11737_n14973.n121 4.5005
R13618 a_n11737_n14973.n64 a_n11737_n14973.n223 4.5005
R13619 a_n11737_n14973.n72 a_n11737_n14973.n71 2.21666
R13620 a_n11737_n14973.n70 a_n11737_n14973.n222 4.5005
R13621 a_n11737_n14973.n87 a_n11737_n14973.n86 2.21666
R13622 a_n11737_n14973.n85 a_n11737_n14973.n221 4.5005
R13623 a_n11737_n14973.n2 a_n11737_n14973.n4 2.21666
R13624 a_n11737_n14973.n91 a_n11737_n14973.n90 2.21666
R13625 a_n11737_n14973.n89 a_n11737_n14973.n217 4.5005
R13626 a_n11737_n14973.n216 a_n11737_n14973.n120 4.5005
R13627 a_n11737_n14973.n60 a_n11737_n14973.n172 4.5005
R13628 a_n11737_n14973.n76 a_n11737_n14973.n75 2.21666
R13629 a_n11737_n14973.n74 a_n11737_n14973.n171 4.5005
R13630 a_n11737_n14973.n94 a_n11737_n14973.n93 0.023589
R13631 a_n11737_n14973.n56 a_n11737_n14973.n55 2.21666
R13632 a_n11737_n14973.n183 a_n11737_n14973.n54 4.5005
R13633 a_n11737_n14973.n42 a_n11737_n14973.n180 4.5005
R13634 a_n11737_n14973.n43 a_n11737_n14973.n45 2.21666
R13635 a_n11737_n14973.n53 a_n11737_n14973.n181 4.5005
R13636 a_n11737_n14973.n80 a_n11737_n14973.n78 2.21666
R13637 a_n11737_n14973.n197 a_n11737_n14973.n196 4.5005
R13638 a_n11737_n14973.n191 a_n11737_n14973.n190 4.5005
R13639 a_n11737_n14973.n189 a_n11737_n14973.n133 4.5005
R13640 a_n11737_n14973.n26 a_n11737_n14973.n177 4.5005
R13641 a_n11737_n14973.n29 a_n11737_n14973.n28 2.21666
R13642 a_n11737_n14973.n27 a_n11737_n14973.n176 4.5005
R13643 a_n11737_n14973.n57 a_n11737_n14973.n59 2.21666
R13644 a_n11737_n14973.n203 a_n11737_n14973.n202 4.5005
R13645 a_n11737_n14973.n47 a_n11737_n14973.n49 4.5005
R13646 a_n11737_n14973.n50 a_n11737_n14973.n48 2.21666
R13647 a_n11737_n14973.n17 a_n11737_n14973.n15 2.21666
R13648 a_n11737_n14973.n199 a_n11737_n14973.n16 4.5005
R13649 a_n11737_n14973.n213 a_n11737_n14973.n212 4.5005
R13650 a_n11737_n14973.n132 a_n11737_n14973.n130 4.5005
R13651 a_n11737_n14973.n131 a_n11737_n14973.n211 4.5005
R13652 a_n11737_n14973.n33 a_n11737_n14973.n31 2.21666
R13653 a_n11737_n14973.n30 a_n11737_n14973.n0 0.0743189
R13654 a_n11737_n14973.n303 a_n11737_n14973.n152 4.5005
R13655 a_n11737_n14973.n283 a_n11737_n14973.n280 4.5005
R13656 a_n11737_n14973.n285 a_n11737_n14973.n284 4.5005
R13657 a_n11737_n14973.n286 a_n11737_n14973.n279 4.5005
R13658 a_n11737_n14973.n288 a_n11737_n14973.n287 4.5005
R13659 a_n11737_n14973.n290 a_n11737_n14973.n289 4.5005
R13660 a_n11737_n14973.n295 a_n11737_n14973.n294 4.5005
R13661 a_n11737_n14973.n119 a_n11737_n14973.n296 4.5005
R13662 a_n11737_n14973.n297 a_n11737_n14973.n153 4.5005
R13663 a_n11737_n14973.n299 a_n11737_n14973.n298 4.5005
R13664 a_n11737_n14973.n300 a_n11737_n14973.n101 4.5005
R13665 a_n11737_n14973.n302 a_n11737_n14973.n301 4.5005
R13666 a_n11737_n14973.n306 a_n11737_n14973.n114 4.5005
R13667 a_n11737_n14973.n308 a_n11737_n14973.n307 4.5005
R13668 a_n11737_n14973.n310 a_n11737_n14973.n151 4.5005
R13669 a_n11737_n14973.n312 a_n11737_n14973.n311 4.5005
R13670 a_n11737_n14973.n313 a_n11737_n14973.n150 4.5005
R13671 a_n11737_n14973.n315 a_n11737_n14973.n314 4.5005
R13672 a_n11737_n14973.n317 a_n11737_n14973.n149 4.5005
R13673 a_n11737_n14973.n327 a_n11737_n14973.n326 4.5005
R13674 a_n11737_n14973.n118 a_n11737_n14973.n116 4.5005
R13675 a_n11737_n14973.n117 a_n11737_n14973.n325 4.5005
R13676 a_n11737_n14973.n324 a_n11737_n14973.n321 4.5005
R13677 a_n11737_n14973.n234 a_n11737_n14973.n226 4.5005
R13678 a_n11737_n14973.n112 a_n11737_n14973.n233 4.5005
R13679 a_n11737_n14973.n232 a_n11737_n14973.n111 4.5005
R13680 a_n11737_n14973.n231 a_n11737_n14973.n230 4.5005
R13681 a_n11737_n14973.n274 a_n11737_n14973.n273 4.5005
R13682 a_n11737_n14973.n272 a_n11737_n14973.n227 4.5005
R13683 a_n11737_n14973.n270 a_n11737_n14973.n269 4.5005
R13684 a_n11737_n14973.n268 a_n11737_n14973.n98 4.5005
R13685 a_n11737_n14973.n267 a_n11737_n14973.n100 4.5005
R13686 a_n11737_n14973.n99 a_n11737_n14973.n238 4.5005
R13687 a_n11737_n14973.n266 a_n11737_n14973.n265 4.5005
R13688 a_n11737_n14973.n254 a_n11737_n14973.n253 4.5005
R13689 a_n11737_n14973.n108 a_n11737_n14973.n255 4.5005
R13690 a_n11737_n14973.n256 a_n11737_n14973.n240 4.5005
R13691 a_n11737_n14973.n258 a_n11737_n14973.n257 4.5005
R13692 a_n11737_n14973.n259 a_n11737_n14973.n97 4.5005
R13693 a_n11737_n14973.n261 a_n11737_n14973.n260 4.5005
R13694 a_n11737_n14973.n262 a_n11737_n14973.n239 4.5005
R13695 a_n11737_n14973.n249 a_n11737_n14973.n248 4.5005
R13696 a_n11737_n14973.n247 a_n11737_n14973.n241 4.5005
R13697 a_n11737_n14973.n246 a_n11737_n14973.n245 4.5005
R13698 a_n11737_n14973.n244 a_n11737_n14973.n242 4.5005
R13699 a_n11737_n14973.n366 a_n11737_n14973.n141 4.5005
R13700 a_n11737_n14973.n134 a_n11737_n14973.n135 2.24296
R13701 a_n11737_n14973.n358 a_n11737_n14973.n357 3.83265
R13702 a_n11737_n14973.n351 a_n11737_n14973.n350 3.82765
R13703 a_n11737_n14973.n134 a_n11737_n14973.t16 3.82673
R13704 a_n11737_n14973.n365 a_n11737_n14973.n364 3.78255
R13705 a_n11737_n14973.n138 a_n11737_n14973.t26 3.76633
R13706 a_n11737_n14973.n372 a_n11737_n14973.n371 3.75068
R13707 a_n11737_n14973.n145 a_n11737_n14973.n144 3.75068
R13708 a_n11737_n14973.n368 a_n11737_n14973.n367 3.74975
R13709 a_n11737_n14973.n225 a_n11737_n14973.n147 3.37223
R13710 a_n11737_n14973.n113 a_n11737_n14973.n305 3.02216
R13711 a_n11737_n14973.n221 a_n11737_n14973.n220 2.89625
R13712 a_n11737_n14973.n18 a_n11737_n14973.n198 2.95081
R13713 a_n11737_n14973.n218 a_n11737_n14973.n163 2.88162
R13714 a_n11737_n14973.n196 a_n11737_n14973.n15 2.95081
R13715 a_n11737_n14973.n344 a_n11737_n14973.n343 2.76066
R13716 a_n11737_n14973.n343 a_n11737_n14973.n342 2.57313
R13717 a_n11737_n14973.n69 a_n11737_n14973.n83 2.00991
R13718 a_n11737_n14973.n276 a_n11737_n14973.n275 2.30989
R13719 a_n11737_n14973.n329 a_n11737_n14973.n148 2.30989
R13720 a_n11737_n14973.n305 a_n11737_n14973.n304 2.29659
R13721 a_n11737_n14973.n264 a_n11737_n14973.n263 2.2812
R13722 a_n11737_n14973.n369 a_n11737_n14973.n368 2.24389
R13723 a_n11737_n14973.n204 a_n11737_n14973.n174 2.23529
R13724 a_n11737_n14973.n186 a_n11737_n14973.n179 2.23529
R13725 a_n11737_n14973.n167 a_n11737_n14973.n165 2.23423
R13726 a_n11737_n14973.n159 a_n11737_n14973.n156 2.23423
R13727 a_n11737_n14973.n289 a_n11737_n14973.n277 2.18975
R13728 a_n11737_n14973.n328 a_n11737_n14973.n149 2.18975
R13729 a_n11737_n14973.n275 a_n11737_n14973.n226 2.16725
R13730 a_n11737_n14973.n254 a_n11737_n14973.n148 2.16725
R13731 a_n11737_n14973.n225 a_n11737_n14973.n224 2.11247
R13732 a_n11737_n14973.n190 a_n11737_n14973.n154 2.102
R13733 a_n11737_n14973.n46 a_n11737_n14973.n213 2.102
R13734 a_n11737_n14973.n362 a_n11737_n14973.n361 2.07395
R13735 a_n11737_n14973.n224 a_n11737_n14973.n154 2.07182
R13736 a_n11737_n14973.n214 a_n11737_n14973.n46 2.07182
R13737 a_n11737_n14973.n37 a_n11737_n14973.n66 2.13751
R13738 a_n11737_n14973.n215 a_n11737_n14973.n62 2.13751
R13739 a_n11737_n14973.n361 a_n11737_n14973.n344 1.90955
R13740 a_n11737_n14973.n336 a_n11737_n14973.n332 1.71486
R13741 a_n11737_n14973.n214 a_n11737_n14973.n147 1.50911
R13742 a_n11737_n14973.n224 a_n11737_n14973.n37 1.5005
R13743 a_n11737_n14973.n215 a_n11737_n14973.n214 1.5005
R13744 a_n11737_n14973.n277 a_n11737_n14973.n276 1.5005
R13745 a_n11737_n14973.n329 a_n11737_n14973.n328 1.5005
R13746 a_n11737_n14973.n336 a_n11737_n14973.n335 1.5005
R13747 a_n11737_n14973.n340 a_n11737_n14973.n339 1.5005
R13748 a_n11737_n14973.n361 a_n11737_n14973.n360 1.5005
R13749 a_n11737_n14973.n371 a_n11737_n14973.t13 1.4705
R13750 a_n11737_n14973.n371 a_n11737_n14973.n370 1.4705
R13751 a_n11737_n14973.n364 a_n11737_n14973.t21 1.4705
R13752 a_n11737_n14973.n364 a_n11737_n14973.n363 1.4705
R13753 a_n11737_n14973.n144 a_n11737_n14973.t24 1.4705
R13754 a_n11737_n14973.n144 a_n11737_n14973.n143 1.4705
R13755 a_n11737_n14973.n348 a_n11737_n14973.t20 1.4705
R13756 a_n11737_n14973.n348 a_n11737_n14973.n347 1.4705
R13757 a_n11737_n14973.n354 a_n11737_n14973.t11 1.4705
R13758 a_n11737_n14973.n354 a_n11737_n14973.n353 1.4705
R13759 a_n11737_n14973.n350 a_n11737_n14973.t27 1.4705
R13760 a_n11737_n14973.n350 a_n11737_n14973.n349 1.4705
R13761 a_n11737_n14973.n283 a_n11737_n14973.n282 1.39514
R13762 a_n11737_n14973.n276 a_n11737_n14973.n225 1.39023
R13763 a_n11737_n14973.n330 a_n11737_n14973.n329 1.39023
R13764 a_n11737_n14973.n146 a_n11737_n14973.n145 1.27228
R13765 a_n11737_n14973.n318 a_n11737_n14973.n317 1.26997
R13766 a_n11737_n14973.n291 a_n11737_n14973.n290 1.26997
R13767 a_n11737_n14973.n326 a_n11737_n14973.n320 1.24392
R13768 a_n11737_n14973.n294 a_n11737_n14973.n293 1.24392
R13769 a_n11737_n14973.n253 a_n11737_n14973.n252 1.24204
R13770 a_n11737_n14973.n235 a_n11737_n14973.n234 1.24204
R13771 a_n11737_n14973.n372 a_n11737_n14973.n369 1.20682
R13772 a_n11737_n14973.n250 a_n11737_n14973.n249 1.20414
R13773 a_n11737_n14973.n273 a_n11737_n14973.n237 1.20414
R13774 a_n11737_n14973.n324 a_n11737_n14973.n323 1.14132
R13775 a_n11737_n14973.n135 a_n11737_n14973.n365 1.20835
R13776 a_n11737_n14973.n231 a_n11737_n14973.n228 1.13598
R13777 a_n11737_n14973.n359 a_n11737_n14973.n351 1.13573
R13778 a_n11737_n14973.n338 a_n11737_n14973.n337 0.90675
R13779 a_n11737_n14973.n334 a_n11737_n14973.n333 0.90675
R13780 a_n11737_n14973.n351 a_n11737_n14973.n137 0.939226
R13781 a_n11737_n14973.n295 a_n11737_n14973.n277 0.752
R13782 a_n11737_n14973.n328 a_n11737_n14973.n327 0.752
R13783 a_n11737_n14973.n275 a_n11737_n14973.n274 0.71825
R13784 a_n11737_n14973.n248 a_n11737_n14973.n148 0.71825
R13785 a_n11737_n14973.n319 a_n11737_n14973.n318 0.663658
R13786 a_n11737_n14973.n320 a_n11737_n14973.n319 0.663658
R13787 a_n11737_n14973.n292 a_n11737_n14973.n291 0.663658
R13788 a_n11737_n14973.n293 a_n11737_n14973.n292 0.663658
R13789 a_n11737_n14973.n251 a_n11737_n14973.n250 0.655156
R13790 a_n11737_n14973.n252 a_n11737_n14973.n251 0.655156
R13791 a_n11737_n14973.n237 a_n11737_n14973.n236 0.655156
R13792 a_n11737_n14973.n236 a_n11737_n14973.n235 0.655156
R13793 a_n11737_n14973.n330 a_n11737_n14973.n147 0.603852
R13794 a_n11737_n14973.n365 a_n11737_n14973.n362 0.596867
R13795 a_n11737_n14973.n96 a_n11737_n14973.n95 0.313126
R13796 a_n11737_n14973.n282 a_n11737_n14973.n281 0.432797
R13797 a_n11737_n14973.n308 a_n11737_n14973.n114 0.394842
R13798 a_n11737_n14973.n303 a_n11737_n14973.n302 0.394842
R13799 a_n11737_n14973.n117 a_n11737_n14973.n321 0.381816
R13800 a_n11737_n14973.n298 a_n11737_n14973.n297 0.381816
R13801 a_n11737_n14973.n245 a_n11737_n14973.n244 0.379447
R13802 a_n11737_n14973.n262 a_n11737_n14973.n261 0.379447
R13803 a_n11737_n14973.n257 a_n11737_n14973.n256 0.379447
R13804 a_n11737_n14973.n270 a_n11737_n14973.n98 0.379447
R13805 a_n11737_n14973.n99 a_n11737_n14973.n266 0.379447
R13806 a_n11737_n14973.n230 a_n11737_n14973.n111 0.379447
R13807 a_n11737_n14973.n182 a_n11737_n14973.n52 0.44431
R13808 a_n11737_n14973.n79 a_n11737_n14973.n195 0.44431
R13809 a_n11737_n14973.n58 a_n11737_n14973.n175 0.44431
R13810 a_n11737_n14973.n1 a_n11737_n14973.n210 1.94004
R13811 a_n11737_n14973.n88 a_n11737_n14973.n105 0.44431
R13812 a_n11737_n14973.n94 a_n11737_n14973.n104 1.95665
R13813 a_n11737_n14973.n56 a_n11737_n14973.n181 0.44431
R13814 a_n11737_n14973.n80 a_n11737_n14973.n176 0.44431
R13815 a_n11737_n14973.n59 a_n11737_n14973.n199 0.44431
R13816 a_n11737_n14973.n301 a_n11737_n14973.n152 0.375125
R13817 a_n11737_n14973.n307 a_n11737_n14973.n306 0.375125
R13818 a_n11737_n14973.n194 a_n11737_n14973.n25 0.431935
R13819 a_n11737_n14973.n32 a_n11737_n14973.n209 0.431935
R13820 a_n11737_n14973.n73 a_n11737_n14973.n107 0.431935
R13821 a_n11737_n14973.n77 a_n11737_n14973.n106 0.431935
R13822 a_n11737_n14973.n29 a_n11737_n14973.n177 0.431935
R13823 a_n11737_n14973.n211 a_n11737_n14973.n33 0.431935
R13824 a_n11737_n14973.n299 a_n11737_n14973.n153 0.36275
R13825 a_n11737_n14973.n325 a_n11737_n14973.n324 0.36275
R13826 a_n11737_n14973.n187 a_n11737_n14973.n178 0.3605
R13827 a_n11737_n14973.n205 a_n11737_n14973.n173 0.3605
R13828 a_n11737_n14973.n160 a_n11737_n14973.n155 0.3605
R13829 a_n11737_n14973.n168 a_n11737_n14973.n166 0.3605
R13830 a_n11737_n14973.n38 a_n11737_n14973.n103 0.3605
R13831 a_n11737_n14973.n223 a_n11737_n14973.n72 0.429685
R13832 a_n11737_n14973.n222 a_n11737_n14973.n87 0.429685
R13833 a_n11737_n14973.n217 a_n11737_n14973.n216 0.3605
R13834 a_n11737_n14973.n172 a_n11737_n14973.n76 0.429685
R13835 a_n11737_n14973.n171 a_n11737_n14973.n94 1.93517
R13836 a_n11737_n14973.n232 a_n11737_n14973.n231 0.3605
R13837 a_n11737_n14973.n269 a_n11737_n14973.n268 0.3605
R13838 a_n11737_n14973.n265 a_n11737_n14973.n238 0.3605
R13839 a_n11737_n14973.n260 a_n11737_n14973.n239 0.3605
R13840 a_n11737_n14973.n258 a_n11737_n14973.n240 0.3605
R13841 a_n11737_n14973.n246 a_n11737_n14973.n242 0.3605
R13842 a_n11737_n14973.n362 a_n11737_n14973.n146 0.339591
R13843 a_n11737_n14973.n323 a_n11737_n14973.n322 0.335806
R13844 a_n11737_n14973.n229 a_n11737_n14973.n228 0.33475
R13845 a_n11737_n14973.n339 a_n11737_n14973.n338 0.320048
R13846 a_n11737_n14973.n335 a_n11737_n14973.n334 0.320048
R13847 a_n11737_n14973.n311 a_n11737_n14973.n150 0.302474
R13848 a_n11737_n14973.n286 a_n11737_n14973.n285 0.302474
R13849 a_n11737_n14973.n185 a_n11737_n14973.n184 0.287375
R13850 a_n11737_n14973.n201 a_n11737_n14973.n200 0.287375
R13851 a_n11737_n14973.n158 a_n11737_n14973.n157 0.287375
R13852 a_n11737_n14973.n164 a_n11737_n14973.n102 0.287375
R13853 a_n11737_n14973.n183 a_n11737_n14973.n180 0.287375
R13854 a_n11737_n14973.n47 a_n11737_n14973.n203 0.287375
R13855 a_n11737_n14973.n284 a_n11737_n14973.n279 0.287375
R13856 a_n11737_n14973.n313 a_n11737_n14973.n312 0.287375
R13857 a_n11737_n14973.n343 a_n11737_n14973.n340 0.212426
R13858 a_n11737_n14973.n160 a_n11737_n14973.n159 0.208888
R13859 a_n11737_n14973.n168 a_n11737_n14973.n165 0.208888
R13860 a_n11737_n14973.n187 a_n11737_n14973.n186 0.20887
R13861 a_n11737_n14973.n205 a_n11737_n14973.n204 0.20887
R13862 a_n11737_n14973.n369 a_n11737_n14973.n141 0.208385
R13863 a_n11737_n14973.n305 a_n11737_n14973.n152 0.208099
R13864 a_n11737_n14973.n264 a_n11737_n14973.n239 0.208099
R13865 a_n11737_n14973.n249 a_n11737_n14973.n241 0.147342
R13866 a_n11737_n14973.n261 a_n11737_n14973.n97 0.147342
R13867 a_n11737_n14973.n256 a_n11737_n14973.n108 0.147342
R13868 a_n11737_n14973.n273 a_n11737_n14973.n272 0.147342
R13869 a_n11737_n14973.n100 a_n11737_n14973.n98 0.147342
R13870 a_n11737_n14973.n112 a_n11737_n14973.n111 0.147342
R13871 a_n11737_n14973.n311 a_n11737_n14973.n310 0.147342
R13872 a_n11737_n14973.n315 a_n11737_n14973.n150 0.147342
R13873 a_n11737_n14973.n118 a_n11737_n14973.n117 0.147342
R13874 a_n11737_n14973.n285 a_n11737_n14973.n280 0.147342
R13875 a_n11737_n14973.n287 a_n11737_n14973.n286 0.147342
R13876 a_n11737_n14973.n297 a_n11737_n14973.n119 0.147342
R13877 a_n11737_n14973.n302 a_n11737_n14973.n101 0.147342
R13878 a_n11737_n14973.n139 a_n11737_n14973.n140 1.2061
R13879 a_n11737_n14973.n355 a_n11737_n14973.n139 0.230885
R13880 a_n11737_n14973.n355 a_n11737_n14973.n345 0.14
R13881 a_n11737_n14973.n136 a_n11737_n14973.n137 1.27228
R13882 a_n11737_n14973.t12 a_n11737_n14973.n136 6.50385
R13883 a_n11737_n14973.n184 a_n11737_n14973.n52 0.209185
R13884 a_n11737_n14973.n185 a_n11737_n14973.n44 0.209185
R13885 a_n11737_n14973.n186 a_n11737_n14973.n44 0.825446
R13886 a_n11737_n14973.n12 a_n11737_n14973.n178 0.209185
R13887 a_n11737_n14973.n7 a_n11737_n14973.n12 0.565419
R13888 a_n11737_n14973.n192 a_n11737_n14973.n7 0.834884
R13889 a_n11737_n14973.n193 a_n11737_n14973.n192 0.14
R13890 a_n11737_n14973.n194 a_n11737_n14973.n193 0.14
R13891 a_n11737_n14973.n195 a_n11737_n14973.n25 0.209185
R13892 a_n11737_n14973.n198 a_n11737_n14973.n79 0.209185
R13893 a_n11737_n14973.n18 a_n11737_n14973.n175 0.209185
R13894 a_n11737_n14973.n201 a_n11737_n14973.n58 0.209185
R13895 a_n11737_n14973.n200 a_n11737_n14973.n51 0.209185
R13896 a_n11737_n14973.n204 a_n11737_n14973.n51 0.825446
R13897 a_n11737_n14973.n14 a_n11737_n14973.n173 0.209185
R13898 a_n11737_n14973.n10 a_n11737_n14973.n14 0.565419
R13899 a_n11737_n14973.n207 a_n11737_n14973.n10 0.834884
R13900 a_n11737_n14973.n208 a_n11737_n14973.n207 0.14
R13901 a_n11737_n14973.n209 a_n11737_n14973.n208 0.14
R13902 a_n11737_n14973.n210 a_n11737_n14973.n32 0.209185
R13903 a_n11737_n14973.n157 a_n11737_n14973.n84 0.209185
R13904 a_n11737_n14973.n158 a_n11737_n14973.n41 0.209185
R13905 a_n11737_n14973.n159 a_n11737_n14973.n41 0.825427
R13906 a_n11737_n14973.n21 a_n11737_n14973.n155 0.209185
R13907 a_n11737_n14973.n162 a_n11737_n14973.n21 0.429685
R13908 a_n11737_n14973.n162 a_n11737_n14973.n129 0.208907
R13909 a_n11737_n14973.n67 a_n11737_n14973.n129 0.836657
R13910 a_n11737_n14973.n67 a_n11737_n14973.n107 0.209185
R13911 a_n11737_n14973.n73 a_n11737_n14973.n105 0.209185
R13912 a_n11737_n14973.n88 a_n11737_n14973.n163 0.209185
R13913 a_n11737_n14973.n218 a_n11737_n14973.n3 0.209185
R13914 a_n11737_n14973.n3 a_n11737_n14973.n92 0.513496
R13915 a_n11737_n14973.n92 a_n11737_n14973.n102 0.209185
R13916 a_n11737_n14973.n36 a_n11737_n14973.n164 0.209185
R13917 a_n11737_n14973.n36 a_n11737_n14973.n165 0.825427
R13918 a_n11737_n14973.n24 a_n11737_n14973.n166 0.209185
R13919 a_n11737_n14973.n170 a_n11737_n14973.n24 0.429685
R13920 a_n11737_n14973.n170 a_n11737_n14973.n126 0.208907
R13921 a_n11737_n14973.n63 a_n11737_n14973.n126 0.836657
R13922 a_n11737_n14973.n63 a_n11737_n14973.n106 0.209185
R13923 a_n11737_n14973.n77 a_n11737_n14973.n104 0.209185
R13924 a_n11737_n14973.n83 a_n11737_n14973.n103 0.209185
R13925 a_n11737_n14973.n39 a_n11737_n14973.n38 0.209137
R13926 a_n11737_n14973.n39 a_n11737_n14973.n37 0.886485
R13927 a_n11737_n14973.n223 a_n11737_n14973.n66 0.209113
R13928 a_n11737_n14973.n222 a_n11737_n14973.n72 0.209185
R13929 a_n11737_n14973.n221 a_n11737_n14973.n87 0.209185
R13930 a_n11737_n14973.n220 a_n11737_n14973.n4 0.209185
R13931 a_n11737_n14973.n91 a_n11737_n14973.n4 0.498871
R13932 a_n11737_n14973.n217 a_n11737_n14973.n91 0.209185
R13933 a_n11737_n14973.n216 a_n11737_n14973.n35 0.209137
R13934 a_n11737_n14973.n215 a_n11737_n14973.n35 0.886485
R13935 a_n11737_n14973.n172 a_n11737_n14973.n62 0.209113
R13936 a_n11737_n14973.n171 a_n11737_n14973.n76 0.209185
R13937 a_n11737_n14973.n56 a_n11737_n14973.n183 0.209185
R13938 a_n11737_n14973.n45 a_n11737_n14973.n180 0.209185
R13939 a_n11737_n14973.n154 a_n11737_n14973.n45 0.908935
R13940 a_n11737_n14973.n190 a_n11737_n14973.n189 0.14
R13941 a_n11737_n14973.n189 a_n11737_n14973.n177 0.14
R13942 a_n11737_n14973.n29 a_n11737_n14973.n176 0.209185
R13943 a_n11737_n14973.n196 a_n11737_n14973.n80 0.209185
R13944 a_n11737_n14973.n199 a_n11737_n14973.n15 0.209185
R13945 a_n11737_n14973.n203 a_n11737_n14973.n59 0.209185
R13946 a_n11737_n14973.n48 a_n11737_n14973.n47 0.209185
R13947 a_n11737_n14973.n48 a_n11737_n14973.n46 0.908935
R13948 a_n11737_n14973.n213 a_n11737_n14973.n130 0.14
R13949 a_n11737_n14973.n211 a_n11737_n14973.n130 0.14
R13950 a_n11737_n14973.n33 a_n11737_n14973.n0 1.54288
R13951 a_n11737_n14973.n284 a_n11737_n14973.n283 0.14
R13952 a_n11737_n14973.n288 a_n11737_n14973.n279 0.14
R13953 a_n11737_n14973.n289 a_n11737_n14973.n288 0.14
R13954 a_n11737_n14973.n296 a_n11737_n14973.n295 0.14
R13955 a_n11737_n14973.n296 a_n11737_n14973.n153 0.14
R13956 a_n11737_n14973.n300 a_n11737_n14973.n299 0.14
R13957 a_n11737_n14973.n301 a_n11737_n14973.n300 0.14
R13958 a_n11737_n14973.n306 a_n11737_n14973.n113 0.208168
R13959 a_n11737_n14973.n307 a_n11737_n14973.n151 0.14
R13960 a_n11737_n14973.n312 a_n11737_n14973.n151 0.14
R13961 a_n11737_n14973.n314 a_n11737_n14973.n313 0.14
R13962 a_n11737_n14973.n314 a_n11737_n14973.n149 0.14
R13963 a_n11737_n14973.n327 a_n11737_n14973.n116 0.14
R13964 a_n11737_n14973.n325 a_n11737_n14973.n116 0.14
R13965 a_n11737_n14973.n233 a_n11737_n14973.n232 0.14
R13966 a_n11737_n14973.n233 a_n11737_n14973.n226 0.14
R13967 a_n11737_n14973.n274 a_n11737_n14973.n227 0.14
R13968 a_n11737_n14973.n269 a_n11737_n14973.n227 0.14
R13969 a_n11737_n14973.n268 a_n11737_n14973.n267 0.14
R13970 a_n11737_n14973.n267 a_n11737_n14973.n238 0.14
R13971 a_n11737_n14973.n265 a_n11737_n14973.n110 0.208168
R13972 a_n11737_n14973.n110 a_n11737_n14973.n264 3.03679
R13973 a_n11737_n14973.n260 a_n11737_n14973.n259 0.14
R13974 a_n11737_n14973.n259 a_n11737_n14973.n258 0.14
R13975 a_n11737_n14973.n255 a_n11737_n14973.n240 0.14
R13976 a_n11737_n14973.n255 a_n11737_n14973.n254 0.14
R13977 a_n11737_n14973.n248 a_n11737_n14973.n247 0.14
R13978 a_n11737_n14973.n247 a_n11737_n14973.n246 0.14
R13979 a_n11737_n14973.n96 a_n11737_n14973.n242 1.12911
R13980 a_n11737_n14973.n141 a_n11737_n14973.n135 0.230894
R13981 a_n11737_n14973.n366 a_n11737_n14973.n134 0.138586
R13982 a_n11737_n14973.n356 a_n11737_n14973.n138 0.137318
R13983 a_n11737_n14973.n230 a_n11737_n14973.n229 0.128395
R13984 a_n11737_n14973.n322 a_n11737_n14973.n321 0.128395
R13985 a_n11737_n14973.n245 a_n11737_n14973.n243 0.118921
R13986 a_n11737_n14973.n263 a_n11737_n14973.n262 0.118921
R13987 a_n11737_n14973.n271 a_n11737_n14973.n270 0.118921
R13988 a_n11737_n14973.n317 a_n11737_n14973.n316 0.114184
R13989 a_n11737_n14973.n290 a_n11737_n14973.n278 0.114184
R13990 a_n11737_n14973.n309 a_n11737_n14973.n308 0.113
R13991 a_n11737_n14973.n358 a_n11737_n14973.n356 0.110782
R13992 a_n11737_n14973.n368 a_n11737_n14973.n366 0.109514
R13993 a_n11737_n14973.n13 a_n11737_n14973.n206 0.109179
R13994 a_n11737_n14973.n11 a_n11737_n14973.n188 0.109179
R13995 a_n11737_n14973.n57 a_n11737_n14973.n16 0.107155
R13996 a_n11737_n14973.n78 a_n11737_n14973.n27 0.107155
R13997 a_n11737_n14973.n55 a_n11737_n14973.n53 0.107155
R13998 a_n11737_n14973.n340 a_n11737_n14973.n336 0.105095
R13999 a_n11737_n14973.n131 a_n11737_n14973.n31 0.103632
R14000 a_n11737_n14973.n28 a_n11737_n14973.n26 0.103632
R14001 a_n11737_n14973.n304 a_n11737_n14973.n303 0.103526
R14002 a_n11737_n14973.n22 a_n11737_n14973.n169 0.102991
R14003 a_n11737_n14973.n124 a_n11737_n14973.n23 0.102991
R14004 a_n11737_n14973.n19 a_n11737_n14973.n161 0.102991
R14005 a_n11737_n14973.n127 a_n11737_n14973.n20 0.102991
R14006 a_n11737_n14973.n360 a_n11737_n14973.n359 0.0995
R14007 a_n11737_n14973.n75 a_n11737_n14973.n60 0.0933826
R14008 a_n11737_n14973.n71 a_n11737_n14973.n64 0.0933826
R14009 a_n11737_n14973.n93 a_n11737_n14973.n74 0.092742
R14010 a_n11737_n14973.n90 a_n11737_n14973.n2 0.092742
R14011 a_n11737_n14973.n86 a_n11737_n14973.n70 0.092742
R14012 a_n11737_n14973.n82 a_n11737_n14973.n68 0.092742
R14013 a_n11737_n14973.n202 a_n11737_n14973.n49 0.0821726
R14014 a_n11737_n14973.n42 a_n11737_n14973.n54 0.0821726
R14015 a_n11737_n14973.n120 a_n11737_n14973.n89 0.0821726
R14016 a_n11737_n14973.n121 a_n11737_n14973.n81 0.0821726
R14017 a_n11737_n14973.n128 a_n11737_n14973.n127 0.0427776
R14018 a_n11737_n14973.n125 a_n11737_n14973.n124 0.0427776
R14019 a_n11737_n14973.n360 a_n11737_n14973.n345 0.041
R14020 a_n11737_n14973.n132 a_n11737_n14973.n131 0.0402153
R14021 a_n11737_n14973.n26 a_n11737_n14973.n133 0.0402153
R14022 a_n11737_n14973.n53 a_n11737_n14973.n122 0.0402153
R14023 a_n11737_n14973.n191 a_n11737_n14973.n133 0.0402153
R14024 a_n11737_n14973.n212 a_n11737_n14973.n132 0.0402153
R14025 a_n11737_n14973.n310 a_n11737_n14973.n309 0.0348421
R14026 a_n11737_n14973.n281 a_n11737_n14973.n280 0.0348421
R14027 a_n11737_n14973.n206 a_n11737_n14973.n174 0.0344623
R14028 a_n11737_n14973.n188 a_n11737_n14973.n179 0.0344623
R14029 a_n11737_n14973.n316 a_n11737_n14973.n315 0.0336579
R14030 a_n11737_n14973.n287 a_n11737_n14973.n278 0.0336579
R14031 a_n11737_n14973.n169 a_n11737_n14973.n167 0.0325285
R14032 a_n11737_n14973.n161 a_n11737_n14973.n156 0.0325285
R14033 a_n11737_n14973.n243 a_n11737_n14973.n241 0.0289211
R14034 a_n11737_n14973.n272 a_n11737_n14973.n271 0.0289211
R14035 a_n11737_n14973.n244 a_n11737_n14973.n95 0.166289
R14036 a_n11737_n14973.n115 a_n11737_n14973.n114 0.156816
R14037 a_n11737_n14973.n266 a_n11737_n14973.n109 0.156816
R14038 a_n11737_n14973.n9 a_n11737_n14973.n8 0.154009
R14039 a_n11737_n14973.n6 a_n11737_n14973.n5 0.154009
R14040 a_n11737_n14973.n294 a_n11737_n14973.n119 0.147342
R14041 a_n11737_n14973.n326 a_n11737_n14973.n118 0.147342
R14042 a_n11737_n14973.n234 a_n11737_n14973.n112 0.147342
R14043 a_n11737_n14973.n253 a_n11737_n14973.n108 0.147342
R14044 a_n11737_n14973.n298 a_n11737_n14973.n101 0.147342
R14045 a_n11737_n14973.n100 a_n11737_n14973.n99 0.147342
R14046 a_n11737_n14973.n257 a_n11737_n14973.n97 0.147342
R14047 a_n11737_n14973.n90 a_n11737_n14973.n89 0.0943434
R14048 a_n11737_n14973.n82 a_n11737_n14973.n81 0.0943434
R14049 a_n11737_n14973.n75 a_n11737_n14973.n74 0.0901797
R14050 a_n11737_n14973.n71 a_n11737_n14973.n70 0.0901797
R14051 a_n11737_n14973.n8 a_n11737_n14973.n13 0.0847264
R14052 a_n11737_n14973.n5 a_n11737_n14973.n11 0.0847264
R14053 a_n11737_n14973.n86 a_n11737_n14973.n85 0.0799306
R14054 a_n11737_n14973.n197 a_n11737_n14973.n78 0.0799306
R14055 a_n11737_n14973.n65 a_n11737_n14973.n64 0.0799306
R14056 a_n11737_n14973.n61 a_n11737_n14973.n60 0.0799306
R14057 a_n11737_n14973.n202 a_n11737_n14973.n57 0.0799306
R14058 a_n11737_n14973.n55 a_n11737_n14973.n54 0.0799306
R14059 a_n11737_n14973.n50 a_n11737_n14973.n49 0.0799306
R14060 a_n11737_n14973.n43 a_n11737_n14973.n42 0.0799306
R14061 a_n11737_n14973.n121 a_n11737_n14973.n40 0.0799306
R14062 a_n11737_n14973.n120 a_n11737_n14973.n34 0.0799306
R14063 a_n11737_n14973.n31 a_n11737_n14973.n30 0.0799306
R14064 a_n11737_n14973.n28 a_n11737_n14973.n27 0.0799306
R14065 a_n11737_n14973.n23 a_n11737_n14973.n22 0.0799306
R14066 a_n11737_n14973.n20 a_n11737_n14973.n19 0.0799306
R14067 a_n11737_n14973.n17 a_n11737_n14973.n16 0.0799306
R14068 a_n11737_n14973.n219 a_n11737_n14973.n2 0.0799306
R14069 a_n11737_n14973.n1 a_n11737_n14973.t107 8.08727
C0 a_n965_n16909# a_n1533_n16909# 0.018349f
C1 a_n2631_n17634# a_n2101_n16909# 0.017843f
C2 a_n1533_n16323# a_n965_n16909# 0.018349f
C3 a_n2101_n16323# a_n1533_n16323# 0.017228f
C4 a_n2631_n16323# a_n2631_n17634# 0.012404f
C5 AVDD IREF 0.25376p
C6 a_n1533_n15598# a_n965_n15598# 0.017228f
C7 a_n2631_n16323# a_n2101_n16323# 0.017843f
C8 a_n2101_n15598# a_n1533_n15598# 0.017228f
C9 a_n1533_n17634# AVDD 0.04859f
C10 IREF VP 0.039954f
C11 AVDD VN 70.0646f
C12 a_n2101_n17634# AVDD 0.030666f
C13 a_n2631_n16323# a_n2101_n15598# 0.017843f
C14 a_n1533_n16909# AVDD 0.016884f
C15 a_n2101_n16909# AVDD 0.016856f
C16 VP VN 55.8707f
C17 a_n2631_n17634# AVDD 0.378896f
C18 a_n965_n16909# AVDD 0.328969f
C19 a_n1533_n16323# AVDD 0.016884f
C20 a_n2101_n16323# AVDD 0.016856f
C21 a_n965_n15598# AVDD 0.165281f
C22 a_n1533_n15598# AVDD 0.030148f
C23 a_n2101_n15598# AVDD 0.030305f
C24 a_n2631_n16323# AVDD 0.378914f
C25 a_n6661_n21443# a_n6139_n21443# 0.017917f
C26 a_n6661_n21443# a_n6139_n20820# 0.017917f
C27 a_n5579_n20820# a_n6139_n20820# 0.017917f
C28 AVDD VP 63.8974f
C29 a_n6139_n20267# a_n5579_n20820# 0.017917f
C30 IREF VN 0.05459f
C31 AVDD VOUT 41.1792f
C32 a_n2101_n17634# a_n1533_n17634# 0.017228f
C33 a_n2101_n16909# a_n1533_n16909# 0.017228f
C34 a_n2631_n17634# a_n2101_n17634# 0.017843f
.ends

