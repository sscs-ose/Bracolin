** sch_path:
*+ /home/gf180/Documents/gf180/gf180_work/PICO_contest/tracking_switches/xschem/on_resistance.sch
**.subckt on_resistance
XM2 Vd Vg GND GND nfet_03v3 L=0.28u W=0.35u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
VDD4 Vg GND 3.3
.save i(vdd4)
VDD1 Vd GND 3.3
.save i(vdd1)
**** begin user architecture code



*Parameters

.options TEMP = 50.0
.lib /home/gf180/Documents/gf180/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.include /home/gf180/Documents/gf180/pdk/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/gf180/Documents/gf180/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/gf180/Documents/gf180/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice mimcap_statistical

*Data to save
.save all


* Simulation
.control

dc VDD4 0 3.3 0.01
plot -i(VDD1)

reset
unset filetype
op
save all
write on_resistance_tb.raw


.endc
.end


**** end user architecture code
**.ends
.GLOBAL GND
.end
