** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_nfets.sch
.subckt FC_nfets S1 S2 D1 D2 G1 G2 B
*.PININFO S1:B S2:B D1:B D2:B G1:B G2:B B:B
M1[1] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[2] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[3] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[4] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[5] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[6] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[7] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[8] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[9] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[10] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[11] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[12] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[13] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[14] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[15] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[16] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[17] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[18] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[1] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[2] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[3] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[4] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[5] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[6] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[7] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[8] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[9] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[10] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[11] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[12] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[13] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[14] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[15] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[16] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[17] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[18] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M3[1] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[2] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[3] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[4] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[5] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[6] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[7] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[8] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[9] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[10] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[11] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[12] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[13] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[14] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[15] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[16] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[17] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[18] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[19] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[20] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[21] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[22] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[23] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[24] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[25] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[26] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[27] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[28] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[29] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[30] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
.ends
.end
