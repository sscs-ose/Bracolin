* Extracted by KLayout with GF180MCU LVS runset on : 01/12/2023 19:06

.SUBCKT FC_net VB2 VB3 VOUT AVDD VP VB4 VN VB1 AVSS
M$1 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$4 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$5 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$6 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$7 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$8 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$9 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$10 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$11 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$12 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$13 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$14 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$15 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$16 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$17 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$18 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$19 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$20 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$21 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$22 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$23 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$24 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$25 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$26 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$27 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$28 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$29 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$30 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$31 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$32 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$33 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$34 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$35 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$36 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$37 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$38 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$39 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$40 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$41 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$42 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$43 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$44 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$45 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$46 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$47 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$48 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$49 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$50 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$51 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$52 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$53 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$54 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$55 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$56 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$57 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$58 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$59 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$60 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$61 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$62 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$63 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$64 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$65 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$66 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$67 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$68 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$69 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$70 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$71 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$72 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$73 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$74 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$75 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$76 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$77 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$78 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$79 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$80 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$81 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$82 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$83 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$84 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$85 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$86 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$87 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$88 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$89 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$90 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$91 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$92 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$93 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$94 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$95 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$96 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$97 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$98 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$99 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$100 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$101 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$102 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$103 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$104 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$105 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$106 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$107 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$108 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$109 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$110 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$111 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$112 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$113 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$114 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$115 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$116 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$117 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$118 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$119 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$120 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$121 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$122 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$123 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$124 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$125 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$126 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$127 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$128 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$129 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$130 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$131 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$132 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$133 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$134 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$135 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$136 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$137 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$138 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$139 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$140 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$141 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$142 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$143 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$144 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$145 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$146 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$147 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$148 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$149 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$150 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$151 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$152 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$153 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$154 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$155 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$156 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$157 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$158 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$159 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$160 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$161 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$162 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$163 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$164 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$165 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$166 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$167 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$168 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$169 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$170 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$171 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$172 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$173 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$174 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$175 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$176 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$177 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$178 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$179 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$180 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$181 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$182 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$183 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$184 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$185 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$186 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$187 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$188 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$189 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$190 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$191 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$192 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$193 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$194 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$195 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$196 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$197 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$198 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$199 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$200 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$201 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$202 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$203 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$204 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$205 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$206 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$207 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$208 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$209 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$210 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$211 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$212 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$213 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$214 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$215 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$216 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$217 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$218 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$219 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$220 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$221 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$222 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$223 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$224 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$225 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$226 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$227 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$228 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$229 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$230 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$231 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$232 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$233 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$234 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$235 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$236 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$237 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$238 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$239 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$240 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$241 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$242 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$243 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$244 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$245 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$246 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$247 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$248 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$249 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$250 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$251 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$252 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$253 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$254 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$255 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$256 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$257 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$258 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$259 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$260 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$261 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$262 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$263 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$264 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$265 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$266 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$267 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$268 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$269 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$270 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$271 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$272 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$273 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$274 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$275 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$276 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$277 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$278 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$279 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$280 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$281 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$282 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$283 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$284 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$285 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$286 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$287 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$288 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$289 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$290 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$291 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$292 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$293 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$294 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$295 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$296 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$297 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$298 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$299 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$300 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$301 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$302 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$303 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$304 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$305 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$306 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$307 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$308 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$309 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$310 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$311 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$312 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$313 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$314 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$315 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$316 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$317 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$318 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$319 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$320 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$321 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$322 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$323 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$324 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$325 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$326 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$327 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$328 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$329 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$330 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$331 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$332 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$333 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$334 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$335 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$336 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$337 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$338 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$339 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$340 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$341 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$342 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$343 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$344 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$345 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$346 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$347 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$348 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$349 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$350 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$351 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$352 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$353 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$354 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$355 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$356 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$357 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$358 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$359 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$360 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$361 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$362 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$363 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$364 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$365 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$366 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$367 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$368 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$369 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$370 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$371 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$372 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$373 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$374 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$375 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$376 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$377 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$378 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$379 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$380 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$381 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$382 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$383 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$384 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$385 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$386 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$387 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$388 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$389 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$390 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$391 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$392 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$393 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$394 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$395 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$396 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$397 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$398 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$399 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$400 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$401 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$402 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$403 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$404 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$405 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$406 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$407 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$408 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$409 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$410 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$411 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$412 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$413 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$414 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$415 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$416 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$417 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$418 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$419 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$420 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$421 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$422 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$423 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$424 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$425 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$426 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$427 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$428 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$429 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$430 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$431 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$432 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$433 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$434 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$435 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$436 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$437 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$438 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$439 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$440 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$441 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$442 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$443 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$444 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$445 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$446 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$447 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$448 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$449 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$450 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$451 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$452 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$453 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$454 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$455 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$456 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$457 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$458 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$459 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$460 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$461 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$462 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$463 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$464 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$465 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$466 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$467 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$468 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$469 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$470 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$471 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$472 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$473 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$474 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$475 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$476 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$477 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$478 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$479 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$480 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$481 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$482 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$483 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$484 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$485 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$486 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$487 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$488 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$489 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$490 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$491 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$492 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$493 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$494 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$495 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$496 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$497 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$498 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$499 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$500 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$501 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$502 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$503 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$504 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$505 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$506 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$507 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$508 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$509 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$510 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$511 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$512 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$513 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$514 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$515 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$516 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$517 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$518 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$519 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$520 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$521 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$522 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$523 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$524 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$525 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$526 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$527 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$528 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$529 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$530 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$531 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$532 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$533 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$534 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$535 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$536 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$537 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$538 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$539 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$540 \$179 VN \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$541 \$14 VN \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$542 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$543 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$544 \$179 VP \$13 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$545 \$13 VP \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$546 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$547 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$548 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$549 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$550 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$551 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$552 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$553 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$554 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$555 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$556 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$557 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$558 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$559 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$560 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$561 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$562 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$563 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$564 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$565 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$566 \$174 VB4 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$567 VOUT VB4 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$568 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$569 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$570 \$180 VB4 \$98 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$571 \$98 VB4 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$572 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$573 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$574 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$575 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$576 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$577 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$578 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$579 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$580 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$581 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$582 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$583 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$584 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$585 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$586 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$587 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$588 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$589 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$590 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$591 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$592 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$593 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$594 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$595 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$596 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$597 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$598 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$599 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$600 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$601 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$602 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$603 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$604 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$605 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$606 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$607 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$608 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$609 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$610 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$611 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$612 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$613 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$614 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$615 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$616 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$617 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$618 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$619 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$620 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$621 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$622 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$623 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$624 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$625 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$626 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$627 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$628 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$629 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$630 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$631 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$632 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$633 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$634 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$635 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$636 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$637 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$638 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$639 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$640 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$641 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$642 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$643 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$644 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$645 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$646 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$647 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$648 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$649 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$650 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$651 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$652 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$653 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$654 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$655 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$656 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$657 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$658 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$659 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$660 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$661 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$662 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$663 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$664 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$665 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$666 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$667 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$668 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$669 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$670 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$671 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$672 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$673 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$674 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$675 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$676 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$677 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$678 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$679 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$680 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$681 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$682 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$683 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$684 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$685 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$686 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$687 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$688 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$689 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$690 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$691 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$692 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$693 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$694 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$695 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$696 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$697 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$698 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$699 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$700 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$701 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$702 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$703 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$704 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$705 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$706 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$707 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$708 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$709 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$710 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$711 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$712 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$713 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$714 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$715 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$716 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$717 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$718 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$719 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$720 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$721 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$722 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$723 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$724 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$725 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$726 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$727 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$728 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$729 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$730 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$731 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$732 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$733 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$734 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$735 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$736 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$737 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$738 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$739 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$740 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$741 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$742 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$743 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$744 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$745 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$746 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$747 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$748 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$749 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$750 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$751 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$752 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$753 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$754 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$755 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$756 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$757 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$758 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$759 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$760 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$761 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$762 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$763 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$764 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$765 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$766 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$767 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$768 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$769 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$770 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$771 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$772 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$773 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$774 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$775 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$776 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$777 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$778 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$779 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$780 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$781 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$782 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$783 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$784 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$785 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$786 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$787 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$788 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$789 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$790 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$791 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$792 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$793 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$794 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$795 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$796 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$797 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$798 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$799 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$800 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$801 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$802 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$803 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$804 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$805 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$806 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$807 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$808 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$809 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$810 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$811 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$812 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$813 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$814 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$815 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$816 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$817 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$818 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$819 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$820 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$821 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$822 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$823 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$824 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$825 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$826 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$827 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$828 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$829 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$830 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$831 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$832 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$833 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$834 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$835 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$836 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$837 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$838 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$839 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$840 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$841 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$842 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$843 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$844 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$845 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$846 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$847 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$848 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$849 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$850 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$851 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$852 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$853 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$854 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$855 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$856 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$857 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$858 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$859 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$860 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$861 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$862 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$863 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$864 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$865 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$866 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$867 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$868 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$869 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$870 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$871 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$872 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$873 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$874 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$875 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$876 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$877 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$878 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$879 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$880 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$881 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$882 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$883 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$884 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$885 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$886 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$887 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$888 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$889 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$890 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$891 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$892 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$893 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$894 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$895 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$896 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$897 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$898 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$899 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$900 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$901 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$902 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$903 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$904 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$905 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$906 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$907 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$908 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$909 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$910 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$911 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$912 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$913 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$914 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$915 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$916 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$917 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$918 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$919 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$920 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$921 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$922 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$923 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$924 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$925 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$926 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$927 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$928 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$929 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$930 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$931 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$932 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$933 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$934 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$935 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$936 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$937 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$938 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$939 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$940 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$941 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$942 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$943 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$944 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$945 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$946 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$947 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$948 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$949 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$950 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$951 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$952 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$953 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$954 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$955 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$956 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$957 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$958 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$959 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$960 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$961 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$962 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$963 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$964 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$965 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$966 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$967 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$968 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$969 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$970 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$971 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$972 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$973 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$974 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$975 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$976 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$977 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$978 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$979 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$980 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$981 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$982 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$983 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$984 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$985 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$986 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$987 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$988 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$989 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$990 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$991 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$992 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$993 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$994 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$995 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$996 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$997 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$998 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$999 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1000 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1001 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1002 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1003 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1004 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1005 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1006 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1007 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1008 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1009 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1010 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1011 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1012 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1013 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1014 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1015 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1016 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1017 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1018 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1019 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1020 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1021 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1022 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1023 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1024 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1025 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1026 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1027 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1028 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1029 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1030 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1031 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1032 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1033 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1034 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1035 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1036 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1037 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1038 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1039 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1040 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1041 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1042 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1043 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1044 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1045 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1046 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1047 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1048 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1049 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1050 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1051 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1052 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1053 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1054 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1055 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1056 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1057 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1058 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1059 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1060 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1061 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1062 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1063 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1064 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1065 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1066 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1067 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1068 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1069 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1070 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1071 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1072 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1073 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1074 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1075 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1076 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1077 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1078 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1079 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1080 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1081 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1082 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1083 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1084 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1085 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1086 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1087 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1088 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1089 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1090 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1091 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1092 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1093 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1094 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1095 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1096 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1097 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1098 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1099 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1100 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1101 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1102 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1103 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1104 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1105 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1106 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1107 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1108 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1109 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1110 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1111 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1112 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1113 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1114 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1115 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1116 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1117 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1118 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1119 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1120 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1121 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1122 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1123 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1124 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1125 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1126 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1127 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1128 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1129 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1130 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1131 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1132 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1133 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1134 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1135 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1136 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1137 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1138 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1139 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1140 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1141 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1142 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1143 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1144 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1145 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1146 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1147 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1148 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1149 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1150 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1151 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1152 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1153 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1154 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1155 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1156 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1157 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1158 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1159 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1160 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1161 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1162 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1163 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1164 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1165 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1166 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1167 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1168 AVDD VB1 \$179 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1169 \$179 VB1 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1170 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1171 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1172 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1173 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1174 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1175 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1176 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1177 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1178 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1179 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1180 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1181 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1182 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1183 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1184 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1185 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1186 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1187 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1188 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1189 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1190 AVDD \$98 \$174 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1191 \$174 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1192 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1193 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1194 AVDD \$98 \$180 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1195 \$180 \$98 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1196 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1197 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1198 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1199 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1200 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1201 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1202 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1203 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1204 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1205 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1206 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1207 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1208 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1209 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1210 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1211 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1212 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1213 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1214 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1215 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1216 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1217 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1218 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1219 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1220 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1221 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1222 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1223 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1224 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1225 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1226 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1227 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1228 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1229 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1230 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1231 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1232 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1233 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1234 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1235 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1236 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1237 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1238 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1239 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1240 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1241 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1242 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1243 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1244 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1245 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1246 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1247 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1248 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1249 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1250 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1251 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1252 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1253 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1254 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1255 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1256 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1257 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1258 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1259 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1260 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1261 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1262 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1263 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1264 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1265 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1266 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1267 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1268 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1269 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1270 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1271 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1272 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1273 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1274 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1275 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1276 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1277 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1278 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1279 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1280 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1281 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1282 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1283 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1284 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1285 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1286 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1287 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1288 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1289 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1290 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1291 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1292 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1293 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1294 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1295 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1296 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1297 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1298 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1299 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1300 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1301 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1302 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1303 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1304 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1305 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1306 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1307 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1308 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1309 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1310 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1311 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1312 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1313 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1314 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1315 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1316 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1317 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1318 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1319 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1320 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1321 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1322 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1323 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1324 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1325 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1326 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1327 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1328 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1329 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1330 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1331 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1332 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1333 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1334 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1335 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1336 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1337 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1338 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1339 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1340 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1341 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1342 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1343 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1344 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1345 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1346 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1347 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1348 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1349 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1350 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1351 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1352 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1353 AVSS VB2 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1354 \$14 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1355 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1356 \$13 VB2 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1357 AVSS VB2 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1358 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1359 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1360 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1361 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1362 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1363 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1364 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1365 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1366 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1367 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1368 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1369 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1370 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1371 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1372 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1373 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1374 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1375 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1376 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1377 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1378 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1379 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1380 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1381 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1382 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1383 \$98 VB3 \$13 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1384 \$13 VB3 \$98 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1385 \$98 VB3 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1386 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1387 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1388 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1389 \$14 VB3 VOUT AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1390 VOUT VB3 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1391 \$14 VB3 VOUT AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1392 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1393 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1394 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1395 \$98 VB3 \$13 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1396 \$13 VB3 \$98 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1397 \$98 VB3 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1398 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1399 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1400 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1401 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1402 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1403 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1404 VOUT VB3 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1405 \$14 VB3 VOUT AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1406 VOUT VB3 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1407 \$98 VB3 \$13 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1408 \$13 VB3 \$98 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1409 \$98 VB3 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1410 \$14 VB3 VOUT AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1411 VOUT VB3 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1412 \$14 VB3 VOUT AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1413 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1414 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1415 VOUT VB3 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1416 \$14 VB3 VOUT AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1417 VOUT VB3 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1418 \$98 VB3 \$13 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1419 \$13 VB3 \$98 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1420 \$98 VB3 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1421 \$14 VB3 VOUT AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1422 VOUT VB3 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1423 \$14 VB3 VOUT AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1424 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1425 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1426 \$98 VB3 \$13 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1427 \$13 VB3 \$98 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1428 \$98 VB3 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1429 VOUT VB3 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1430 \$14 VB3 VOUT AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1431 VOUT VB3 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1432 \$13 VB3 \$98 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1433 \$98 VB3 \$13 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1434 \$13 VB3 \$98 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1435 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1436 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1437 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1438 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1439 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1440 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1441 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1442 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1443 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1444 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1445 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1446 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
.ENDS FC_net
