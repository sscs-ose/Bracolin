* Extracted by KLayout with GF180MCU LVS runset on : 05/04/2024 17:26

.SUBCKT Res_Div GND vref_off Vout
R$1 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$2 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$3 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$4 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$5 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$6 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$7 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$8 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$9 \$3 \$4 GND 5000 ppolyf_u_1k L=10U W=2U
R$10 \$4 \$5 GND 5000 ppolyf_u_1k L=10U W=2U
R$11 \$5 \$6 GND 5000 ppolyf_u_1k L=10U W=2U
R$12 \$6 \$7 GND 5000 ppolyf_u_1k L=10U W=2U
R$13 \$7 \$8 GND 5000 ppolyf_u_1k L=10U W=2U
R$14 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$15 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$16 \$3 \$11 GND 5000 ppolyf_u_1k L=10U W=2U
R$17 \$11 \$12 GND 5000 ppolyf_u_1k L=10U W=2U
R$18 \$12 \$13 GND 5000 ppolyf_u_1k L=10U W=2U
R$19 \$13 \$14 GND 5000 ppolyf_u_1k L=10U W=2U
R$20 \$14 vref_off GND 5000 ppolyf_u_1k L=10U W=2U
R$21 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$22 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$23 Vout \$17 GND 5000 ppolyf_u_1k L=10U W=2U
R$24 \$17 \$18 GND 5000 ppolyf_u_1k L=10U W=2U
R$25 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$26 \$18 \$19 GND 5000 ppolyf_u_1k L=10U W=2U
R$27 \$19 vref_off GND 5000 ppolyf_u_1k L=10U W=2U
R$28 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$29 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$30 \$26 \$27 GND 5000 ppolyf_u_1k L=10U W=2U
R$31 \$27 \$28 GND 5000 ppolyf_u_1k L=10U W=2U
R$32 \$28 \$29 GND 5000 ppolyf_u_1k L=10U W=2U
R$33 \$29 \$30 GND 5000 ppolyf_u_1k L=10U W=2U
R$34 \$30 \$8 GND 5000 ppolyf_u_1k L=10U W=2U
R$35 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$36 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$37 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$38 \$26 \$35 GND 5000 ppolyf_u_1k L=10U W=2U
R$39 \$35 \$36 GND 5000 ppolyf_u_1k L=10U W=2U
R$40 \$36 \$37 GND 5000 ppolyf_u_1k L=10U W=2U
R$41 \$37 GND GND 5000 ppolyf_u_1k L=10U W=2U
R$42 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$43 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$44 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$45 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$46 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$47 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$48 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
R$49 GND GND GND 5000 ppolyf_u_1k L=10U W=2U
.ENDS Res_Div
