* NGSPICE file created from PR_nfets.ext - technology: gf180mcuD

.subckt PR_nfets VD2 VG VC VS2 VS1 VD1 VB
X0 VB.t71 VB.t70 VB.t71 VB.t8 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1 a_430_3128# VG.t0 VS2.t0 VB.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2 a_430_1204# VG.t1 VD1.t1 VB.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3 VB.t69 VB.t68 VB.t69 VB.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4 a_1834_46# VG.t2 VC.t3 VB.t0 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5 a_430_46# VG.t3 VD2.t1 VB.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6 VB.t67 VB.t66 VB.t67 VB.t20 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X7 a_1834_1970# VG.t4 VS1.t3 VB.t0 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X8 VD1 VG.t5 a_1834_1970# VB.t2 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X9 VB.t65 VB.t64 VB.t65 VB.t8 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X10 VB.t63 VB.t62 VB.t63 VB.t20 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X11 VB.t61 VB.t60 VB.t61 VB.t15 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X12 VB.t59 VB.t58 VB.t59 VB.t8 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X13 VB.t57 VB.t56 VB.t57 VB.t2 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X14 VC VG.t6 a_430_3128# VB.t1 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X15 VB.t55 VB.t54 VB.t55 VB.t15 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X16 VB.t53 VB.t52 VB.t53 VB.t20 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X17 VB.t51 VB.t50 VB.t51 VB.t0 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X18 VB.t49 VB.t48 VB.t49 VB.t8 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X19 a_430_1970# VG.t7 VD1.t2 VB.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X20 VS1 VG.t8 a_430_1204# VB.t1 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X21 VB.t47 VB.t46 VB.t47 VB.t3 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X22 VB.t45 VB.t44 VB.t45 VB.t0 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X23 VB.t43 VB.t42 VB.t43 VB.t2 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X24 VB.t41 VB.t40 VB.t41 VB.t8 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X25 VB.t39 VB.t38 VB.t39 VB.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X26 VB.t37 VB.t36 VB.t37 VB.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X27 VB.t35 VB.t34 VB.t35 VB.t3 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X28 VB.t33 VB.t32 VB.t33 VB.t20 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X29 VB.t31 VB.t30 VB.t31 VB.t15 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X30 VB.t29 VB.t28 VB.t29 VB.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X31 VC VG.t9 a_430_46# VB.t1 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X32 VB.t27 VB.t26 VB.t27 VB.t20 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X33 VS1 VG.t10 a_430_1970# VB.t1 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X34 VB.t25 VB.t24 VB.t25 VB.t15 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X35 VB.t23 VB.t22 VB.t23 VB.t1 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X36 VB.t21 VB.t19 VB.t21 VB.t20 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X37 VB.t18 VB.t17 VB.t18 VB.t15 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X38 VS2 VG.t11 a_1834_46# VB.t2 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X39 VB.t16 VB.t14 VB.t16 VB.t15 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X40 VB.t13 VB.t12 VB.t13 VB.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X41 VB.t11 VB.t10 VB.t11 VB.t1 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X42 a_1834_3128# VG.t12 VC.t1 VB.t0 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X43 VD2 VG.t13 a_1834_3128# VB.t2 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X44 VD1 VG.t14 a_1834_1204# VB.t2 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X45 VB.t9 VB.t7 VB.t9 VB.t8 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X46 a_1834_1204# VG.t15 VS1.t0 VB.t0 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X47 VB.t6 VB.t4 VB.t6 VB.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
R0 VB.n58 VB.n6 523.342
R1 VB.n61 VB.n5 521.869
R2 VB.n58 VB.n5 519.659
R3 VB.n61 VB.n6 516.342
R4 VB.t2 VB.t8 452.031
R5 VB.t3 VB.t5 452.031
R6 VB.t8 VB.t20 307.954
R7 VB.t0 VB.t2 307.954
R8 VB.t1 VB.t3 307.954
R9 VB.t5 VB.t15 307.954
R10 VB.t20 VB.n5 256.899
R11 VB.t15 VB.n6 256.899
R12 VB.n59 VB.t0 221.066
R13 VB.n60 VB.t1 215.567
R14 VB.n60 VB.n59 27.4963
R15 VB.n20 VB.t40 8.06917
R16 VB.n20 VB.t19 8.06917
R17 VB.n18 VB.t7 8.06917
R18 VB.n18 VB.t66 8.06917
R19 VB.n17 VB.t64 8.06917
R20 VB.n17 VB.t32 8.06917
R21 VB.n13 VB.t70 8.06917
R22 VB.n13 VB.t62 8.06917
R23 VB.n12 VB.t58 8.06917
R24 VB.n12 VB.t52 8.06917
R25 VB.n69 VB.t48 8.06917
R26 VB.n69 VB.t26 8.06917
R27 VB.n53 VB.t34 8.06917
R28 VB.n27 VB.t10 8.06917
R29 VB.n7 VB.t44 8.06917
R30 VB.n23 VB.t42 8.06917
R31 VB.n50 VB.t14 8.06917
R32 VB.n50 VB.t68 8.06917
R33 VB.n48 VB.t60 8.06917
R34 VB.n48 VB.t38 8.06917
R35 VB.n47 VB.t30 8.06917
R36 VB.n47 VB.t12 8.06917
R37 VB.n43 VB.t54 8.06917
R38 VB.n43 VB.t36 8.06917
R39 VB.n42 VB.t17 8.06917
R40 VB.n42 VB.t28 8.06917
R41 VB.n40 VB.t24 8.06917
R42 VB.n40 VB.t4 8.06917
R43 VB.n34 VB.t46 8.06917
R44 VB.n35 VB.t22 8.06917
R45 VB.n64 VB.t50 8.06917
R46 VB.n3 VB.t56 8.06917
R47 VB.n52 VB.t35 3.3605
R48 VB.n56 VB.t11 3.3605
R49 VB.n26 VB.t45 3.3605
R50 VB.n22 VB.t43 3.3605
R51 VB.n38 VB.t47 3.3605
R52 VB.t23 VB.n4 3.3605
R53 VB.n63 VB.t51 3.3605
R54 VB.n67 VB.t57 3.3605
R55 VB.n66 VB.n65 2.1005
R56 VB.n37 VB.n36 2.1005
R57 VB.n25 VB.n24 2.1005
R58 VB.n55 VB.n54 2.1005
R59 VB.t11 VB.n55 1.2605
R60 VB.n55 VB.t35 1.2605
R61 VB.n25 VB.t43 1.2605
R62 VB.t45 VB.n25 1.2605
R63 VB.n37 VB.t23 1.2605
R64 VB.t47 VB.n37 1.2605
R65 VB.t57 VB.n66 1.2605
R66 VB.n66 VB.t51 1.2605
R67 VB.n8 VB.t21 0.918039
R68 VB.n9 VB.t67 0.918039
R69 VB.n10 VB.t33 0.918039
R70 VB.n11 VB.t63 0.918039
R71 VB.n0 VB.t53 0.918039
R72 VB.n2 VB.t27 0.918039
R73 VB.n28 VB.t69 0.918039
R74 VB.n29 VB.t39 0.918039
R75 VB.n30 VB.t13 0.918039
R76 VB.n31 VB.t37 0.918039
R77 VB.n32 VB.t29 0.918039
R78 VB.n33 VB.t6 0.918039
R79 VB.n8 VB.t41 0.91749
R80 VB.n9 VB.t9 0.91749
R81 VB.n10 VB.t65 0.91749
R82 VB.n11 VB.t71 0.91749
R83 VB.n0 VB.t59 0.91749
R84 VB.n2 VB.t49 0.91749
R85 VB.n28 VB.t16 0.91749
R86 VB.n29 VB.t61 0.91749
R87 VB.n30 VB.t31 0.91749
R88 VB.n31 VB.t55 0.91749
R89 VB.n32 VB.t18 0.91749
R90 VB.n33 VB.t25 0.91749
R91 VB.n39 VB.n33 0.582999
R92 VB.n41 VB.n32 0.582999
R93 VB.n44 VB.n31 0.582999
R94 VB.n46 VB.n30 0.582999
R95 VB.n49 VB.n29 0.582999
R96 VB.n51 VB.n28 0.582999
R97 VB.n68 VB.n2 0.582999
R98 VB.n1 VB.n0 0.582999
R99 VB.n14 VB.n11 0.582999
R100 VB.n16 VB.n10 0.582999
R101 VB.n19 VB.n9 0.582999
R102 VB.n21 VB.n8 0.582999
R103 VB.n45 VB.n6 0.0886356
R104 VB.n58 VB.n57 0.0886356
R105 VB.n59 VB.n58 0.0886356
R106 VB.n15 VB.n5 0.0886356
R107 VB.n62 VB.n61 0.0871667
R108 VB.n61 VB.n60 0.0871667
R109 VB.n50 VB.n49 0.0390622
R110 VB.n41 VB.n40 0.0390622
R111 VB.n20 VB.n19 0.0385696
R112 VB.n48 VB.n47 0.0371211
R113 VB.n43 VB.n42 0.0371211
R114 VB.n18 VB.n17 0.0366533
R115 VB.n13 VB.n12 0.0366533
R116 VB.n23 VB.n22 0.0341
R117 VB.n24 VB.n23 0.0341
R118 VB.n24 VB.n7 0.0341
R119 VB.n26 VB.n7 0.0341
R120 VB.n56 VB.n27 0.0341
R121 VB.n54 VB.n27 0.0341
R122 VB.n54 VB.n53 0.0341
R123 VB.n53 VB.n52 0.0341
R124 VB.n39 VB.n38 0.0302339
R125 VB.n46 VB.n45 0.0301981
R126 VB.n68 VB.n67 0.0301505
R127 VB.n52 VB.n51 0.0300328
R128 VB.n22 VB.n21 0.0299989
R129 VB.n16 VB.n15 0.0298187
R130 VB.n67 VB.n3 0.0294988
R131 VB.n65 VB.n3 0.0294988
R132 VB.n65 VB.n64 0.0294988
R133 VB.n64 VB.n63 0.0294988
R134 VB.n35 VB.n4 0.0294988
R135 VB.n36 VB.n35 0.0294988
R136 VB.n36 VB.n34 0.0294988
R137 VB.n38 VB.n34 0.0294988
R138 VB VB.n1 0.0289244
R139 VB.n45 VB.n44 0.0203634
R140 VB.n15 VB.n14 0.0201097
R141 VB.n57 VB.n56 0.01994
R142 VB.n51 VB.n50 0.0196517
R143 VB.n49 VB.n48 0.0196517
R144 VB.n47 VB.n46 0.0196517
R145 VB.n44 VB.n43 0.0196517
R146 VB.n42 VB.n41 0.0196517
R147 VB.n40 VB.n39 0.0196517
R148 VB.n21 VB.n20 0.019407
R149 VB.n19 VB.n18 0.019407
R150 VB.n17 VB.n16 0.019407
R151 VB.n14 VB.n13 0.019407
R152 VB.n12 VB.n1 0.019407
R153 VB.n69 VB.n68 0.019407
R154 VB.n63 VB.n62 0.0183136
R155 VB.n57 VB.n26 0.01514
R156 VB.n62 VB.n4 0.0120995
R157 VB VB.n69 0.0101451
R158 VG.n1 VG.t13 8.40342
R159 VG.n8 VG.t5 8.40342
R160 VG.n16 VG.t14 8.40342
R161 VG.n24 VG.t11 8.40342
R162 VG.n1 VG.t12 8.32322
R163 VG.n8 VG.t4 8.32322
R164 VG.n16 VG.t15 8.32322
R165 VG.n24 VG.t2 8.32322
R166 VG.n28 VG.t3 8.14051
R167 VG.n5 VG.t0 8.14051
R168 VG.n12 VG.t7 8.14051
R169 VG.n20 VG.t1 8.14051
R170 VG.n26 VG.t9 8.06917
R171 VG.n3 VG.t6 8.06917
R172 VG.n10 VG.t10 8.06917
R173 VG.n18 VG.t8 8.06917
R174 VG.n4 VG.n0 4.5005
R175 VG.n11 VG.n7 4.5005
R176 VG.n19 VG.n15 4.5005
R177 VG.n27 VG.n23 4.5005
R178 VG.n3 VG.n2 2.27692
R179 VG.n10 VG.n9 2.27692
R180 VG.n18 VG.n17 2.27692
R181 VG.n26 VG.n25 2.27692
R182 VG.n6 VG.n5 1.90721
R183 VG.n13 VG.n12 1.90721
R184 VG.n21 VG.n20 1.90721
R185 VG.n29 VG.n28 1.90721
R186 VG.n2 VG.n1 1.72165
R187 VG.n9 VG.n8 1.72165
R188 VG.n17 VG.n16 1.72165
R189 VG.n25 VG.n24 1.72165
R190 VG.n14 VG.n6 1.67138
R191 VG.n22 VG.n21 1.5005
R192 VG.n14 VG.n13 1.5005
R193 VG.n30 VG.n29 1.5005
R194 VG.n5 VG.n4 0.472163
R195 VG.n12 VG.n11 0.472163
R196 VG.n20 VG.n19 0.472163
R197 VG.n22 VG.n14 0.414926
R198 VG VG.n27 0.248
R199 VG VG.n30 0.235838
R200 VG.n2 VG.n0 0.234207
R201 VG.n9 VG.n7 0.234207
R202 VG.n17 VG.n15 0.234207
R203 VG.n25 VG.n23 0.234207
R204 VG.n28 VG 0.224663
R205 VG.n30 VG.n22 0.171682
R206 VG.n4 VG.n3 0.118921
R207 VG.n11 VG.n10 0.118921
R208 VG.n19 VG.n18 0.118921
R209 VG.n27 VG.n26 0.118921
R210 VG.n6 VG.n0 0.0474014
R211 VG.n13 VG.n7 0.0474014
R212 VG.n21 VG.n15 0.0474014
R213 VG.n29 VG.n23 0.0474014
R214 VS2.n1 VS2.t0 11.1022
R215 VS2.n1 VS2 5.50993
R216 VS2 VS2.n0 3.78563
R217 VS2 VS2.n1 0.51665
R218 VD1.n4 VD1.n0 5.28726
R219 VD1.n0 VD1.t2 3.8555
R220 VD1.n3 VD1.n1 3.85313
R221 VD1.n0 VD1.t1 3.68261
R222 VD1 VD1.n2 3.61511
R223 VD1 VD1.n4 2.01431
R224 VD1.n4 VD1.n3 1.54399
R225 VD1.n3 VD1 0.0703684
R226 VC.n4 VC.n1 5.35163
R227 VC.n4 VC.n3 4.49014
R228 VC.n1 VC.t1 4.1605
R229 VC.n3 VC.t3 4.15932
R230 VC.n1 VC.n0 4.15747
R231 VC VC.n2 3.79392
R232 VC VC.n4 0.456321
R233 VC.n3 VC 0.362863
R234 VD2.n1 VD2.n0 10.3339
R235 VD2.n1 VD2 5.95212
R236 VD2 VD2.t1 3.7205
R237 VD2 VD2.n1 0.3893
R238 VS1.n3 VS1.n2 3.84484
R239 VS1.n0 VS1.t3 3.69326
R240 VS1.n3 VS1.n1 3.69326
R241 VS1 VS1.t0 3.61511
R242 VS1 VS1.n4 3.58734
R243 VS1.n0 VS1 0.230237
R244 VS1.n4 VS1.n3 0.188652
R245 VS1.n4 VS1.n0 0.132718
C0 VD2 a_1834_3128# 0.0284f
C1 VG a_430_1970# 0.158107f
C2 a_430_1970# VS1 0.042325f
C3 VD2 a_430_46# 0.029617f
C4 VG a_1834_1970# 0.132223f
C5 VG VS1 1.68829f
C6 a_1834_1970# VS1 0.076822f
C7 VD1 a_430_1970# 0.029136f
C8 VG VC 2.16294f
C9 VG a_1834_46# 0.130866f
C10 VC VS1 0.30855f
C11 a_1834_46# VS1 0.035176f
C12 a_1834_46# VC 0.0284f
C13 VG a_430_3128# 0.157107f
C14 a_430_3128# VC 0.034548f
C15 VS2 VG 2.82601f
C16 a_430_1204# VG 0.158104f
C17 VG VD1 1.07843f
C18 VS2 VS1 1.25935f
C19 a_1834_1970# VD1 0.03168f
C20 a_430_1204# VS1 0.029151f
C21 VD1 VS1 2.76284f
C22 VG a_1834_3128# 0.130866f
C23 a_1834_3128# VS1 0.035176f
C24 VS2 VC 2.53042f
C25 VS2 a_1834_46# 0.029465f
C26 VD1 VC 0.26328f
C27 VG a_430_46# 0.157107f
C28 a_1834_3128# VC 0.0284f
C29 VS2 a_430_3128# 0.0284f
C30 VG a_1834_1204# 0.132223f
C31 VG VD2 4.32433f
C32 a_430_46# VC 0.034548f
C33 a_1834_1204# VS1 0.063642f
C34 VD2 VS1 0.339679f
C35 VD2 VC 2.5807f
C36 VS2 VD1 0.426992f
C37 a_430_1204# VD1 0.042519f
C38 VS2 VD2 2.39841f
C39 VD1 a_1834_1204# 0.045063f
C40 VD1 VD2 0.363029f
.ends

