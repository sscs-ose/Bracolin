* NGSPICE file created from FC_top.ext - technology: gf180mcuD

.subckt FC_top VP VN VOUT IREF AVSS AVDD
X0 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3 a_n11737_n15980# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X7 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X8 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X9 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X10 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X11 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X12 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X13 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X14 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X15 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X16 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X17 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X18 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X19 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X20 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X21 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X22 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X23 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X24 a_n11737_n15980# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X25 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X26 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X27 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X28 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X29 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X30 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X31 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X32 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X33 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X34 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X35 AVDD IREF IREF AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X36 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X37 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X38 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X39 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X40 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X41 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X42 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X43 a_n11737_n15980# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X44 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X45 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X46 AVDD IREF a_n11737_n14973# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X47 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X48 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X49 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X50 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X51 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X52 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X53 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X54 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X55 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X56 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X57 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X58 a_n1533_n15598# a_n11317_n20927# a_n2101_n15598# AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X59 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X60 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X61 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X62 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X63 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X64 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X65 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X66 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X67 AVDD IREF a_n11737_n15980# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X68 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X69 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X70 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X71 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X72 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X73 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X74 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X75 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X76 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X77 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X78 a_n13990_n6451# a_n11737_n15980# a_5396_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X79 a_n11317_n20927# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X80 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X81 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X82 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X83 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X84 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X85 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X86 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X87 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X88 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X89 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X90 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X91 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X92 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X93 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X94 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X95 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X96 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X97 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X98 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X99 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X100 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X101 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X102 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X103 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X104 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X105 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X106 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X107 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X108 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X109 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X110 a_n1533_n16323# a_n11317_n20927# a_n2101_n16323# AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X111 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X112 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X113 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X114 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X115 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X116 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X117 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X118 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X119 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X120 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X121 IREF IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X122 a_n11737_n14973# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X123 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X124 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X125 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X126 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X127 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X128 AVDD IREF a_n11737_n15980# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X129 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X130 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X131 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X132 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X133 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X134 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X135 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X136 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X137 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X138 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X139 a_n2101_n15598# a_n11317_n20927# a_n2631_n16323# AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X140 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X141 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X142 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X143 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X144 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X145 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X146 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X147 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X148 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X149 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X150 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X151 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X152 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X153 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X154 a_n13990_n5465# a_n11737_n15980# VOUT AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X155 a_n13990_n5465# a_n11737_n15980# VOUT AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X156 AVDD IREF a_n11737_n15980# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X157 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X158 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X159 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X160 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X161 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X162 IREF IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X163 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X164 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X165 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X166 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X167 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X168 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X169 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X170 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X171 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X172 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X173 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X174 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X175 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X176 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X177 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X178 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X179 AVDD IREF a_n11737_n14973# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X180 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X181 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X182 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X183 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X184 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X185 AVDD IREF a_n11737_n14973# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X186 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X187 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X188 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X189 a_n2101_n16323# a_n11317_n20927# a_n2631_n16323# AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X190 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X191 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X192 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X193 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X194 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X195 a_n6139_n21443# a_n11737_n15980# a_n6661_n21443# AVSS nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X196 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X197 a_n13990_n5465# a_n11737_n15980# VOUT AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X198 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X199 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X200 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X201 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X202 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X203 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X204 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X205 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X206 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X207 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X208 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X209 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X210 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X211 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X212 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X213 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X214 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X215 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X216 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X217 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X218 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X219 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X220 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X221 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X222 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X223 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X224 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X225 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X226 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X227 a_n1533_n17634# a_n11317_n20927# a_n2101_n17634# AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X228 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X229 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X230 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X231 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X232 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X233 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X234 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X235 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X236 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X237 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X238 a_5396_n6451# a_n11737_n15980# a_n13990_n6451# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X239 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X240 a_5396_n6451# a_n11737_n15980# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X241 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X242 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X243 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X244 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X245 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X246 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X247 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X248 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X249 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X250 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X251 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X252 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X253 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X254 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X255 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X256 AVDD IREF IREF AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X257 AVDD IREF IREF AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X258 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X259 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X260 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X261 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X262 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X263 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X264 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X265 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X266 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X267 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X268 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X269 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X270 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X271 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X272 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X273 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X274 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X275 a_n11737_n14973# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X276 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X277 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X278 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X279 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X280 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X281 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X282 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X283 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X284 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X285 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X286 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X287 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X288 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X289 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X290 a_5396_n6451# a_n11737_n15980# a_n13990_n6451# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X291 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X292 a_5396_n6451# a_n11737_n15980# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X293 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X294 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X295 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X296 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X297 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X298 a_n13990_n6451# a_n11737_n15980# a_5396_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X299 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X300 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X301 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X302 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X303 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X304 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X305 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X306 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X307 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X308 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X309 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X310 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X311 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X312 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X313 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X314 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X315 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X316 a_n2101_n17634# a_n11317_n20927# a_n2631_n17634# AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X317 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X318 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X319 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X320 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X321 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X322 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X323 IREF IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X324 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X325 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X326 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X327 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X328 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X329 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X330 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X331 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X332 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X333 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X334 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X335 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X336 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X337 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X338 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X339 IREF IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X340 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X341 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X342 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X343 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X344 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X345 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X346 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X347 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X348 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X349 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X350 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X351 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X352 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X353 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X354 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X355 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X356 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X357 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X358 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X359 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X360 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X361 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X362 a_n13990_n5465# a_n11737_n15980# VOUT AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X363 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X364 a_n13990_n5465# a_n11737_n15980# VOUT AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X365 a_n6139_n20820# a_n11737_n15980# a_n6661_n21443# AVSS nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X366 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X367 VOUT a_n11737_n15980# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X368 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X369 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X370 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X371 AVDD IREF a_n11737_n14973# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X372 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X373 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X374 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X375 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X376 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X377 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X378 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X379 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X380 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X381 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X382 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X383 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X384 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X385 AVDD IREF IREF AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X386 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X387 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X388 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X389 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X390 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X391 AVDD IREF a_n11737_n15980# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X392 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X393 a_n965_n16909# a_n11317_n20927# a_n1533_n16909# AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X394 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X395 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X396 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X397 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X398 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X399 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X400 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X401 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X402 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X403 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X404 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X405 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X406 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X407 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X408 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X409 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X410 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X411 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X412 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X413 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X414 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X415 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X416 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X417 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X418 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X419 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X420 AVSS a_n11737_n14973# a_n11737_n14973# AVSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X421 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X422 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X423 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X424 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X425 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X426 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X427 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X428 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X429 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X430 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X431 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X432 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X433 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X434 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X435 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X436 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X437 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X438 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X439 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X440 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X441 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X442 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X443 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X444 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X445 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X446 a_n11737_n14973# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X447 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X448 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X449 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X450 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X451 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X452 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X453 a_5396_n6451# a_n11737_n15980# a_n13990_n6451# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X454 AVSS a_n11737_n14973# a_n11317_n20927# AVSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X455 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X456 a_5396_n6451# a_n11737_n15980# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X457 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X458 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X459 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X460 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X461 a_n11737_n14973# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X462 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X463 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X464 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X465 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X466 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X467 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X468 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X469 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X470 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X471 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X472 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X473 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X474 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X475 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X476 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X477 a_n11737_n15980# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X478 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X479 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X480 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X481 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X482 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X483 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X484 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X485 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X486 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X487 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X488 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X489 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X490 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X491 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X492 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X493 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X494 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X495 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X496 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X497 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X498 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X499 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X500 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X501 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X502 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X503 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X504 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X505 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X506 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X507 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X508 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X509 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X510 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X511 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X512 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X513 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X514 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X515 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X516 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X517 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X518 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X519 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X520 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X521 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X522 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X523 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X524 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X525 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X526 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X527 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X528 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X529 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X530 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X531 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X532 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X533 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X534 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X535 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X536 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X537 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X538 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X539 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X540 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X541 IREF IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X542 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X543 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X544 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X545 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X546 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X547 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X548 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X549 a_n13990_n5465# a_n11737_n15980# VOUT AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X550 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X551 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X552 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X553 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X554 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X555 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X556 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X557 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X558 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X559 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X560 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X561 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X562 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X563 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X564 AVDD IREF a_n11737_n14973# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X565 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X566 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X567 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X568 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X569 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X570 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X571 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X572 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X573 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X574 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X575 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X576 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X577 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X578 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X579 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X580 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X581 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X582 VOUT a_n11737_n15980# a_n13990_n5465# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X583 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X584 VOUT a_n11737_n15980# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X585 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X586 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X587 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X588 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X589 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X590 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X591 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X592 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X593 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X594 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X595 AVDD IREF a_n11737_n14973# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X596 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X597 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X598 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X599 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X600 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X601 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X602 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X603 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X604 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X605 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X606 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X607 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X608 AVDD IREF IREF AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X609 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X610 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X611 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X612 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X613 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X614 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X615 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X616 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X617 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X618 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X619 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X620 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X621 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X622 a_5396_n6451# a_n11737_n15980# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X623 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X624 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X625 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X626 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X627 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X628 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X629 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X630 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X631 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X632 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X633 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X634 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X635 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X636 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X637 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X638 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X639 a_n11737_n15980# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X640 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X641 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X642 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X643 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X644 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X645 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X646 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X647 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X648 IREF IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X649 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X650 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X651 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X652 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X653 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X654 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X655 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X656 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X657 a_n11737_n14973# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X658 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X659 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X660 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X661 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X662 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X663 a_n965_n15598# a_n11317_n20927# a_n1533_n15598# AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X664 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X665 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X666 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X667 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X668 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X669 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X670 a_n11737_n15980# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X671 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X672 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X673 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X674 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X675 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X676 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X677 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X678 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X679 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X680 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X681 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X682 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X683 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X684 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X685 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X686 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X687 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X688 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X689 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X690 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X691 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X692 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X693 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X694 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X695 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X696 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X697 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X698 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X699 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X700 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X701 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X702 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X703 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X704 AVDD IREF a_n11737_n15980# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X705 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X706 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X707 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X708 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X709 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X710 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X711 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X712 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X713 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X714 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X715 a_n965_n16909# a_n11317_n20927# a_n1533_n16323# AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X716 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X717 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X718 AVDD IREF a_n11737_n14973# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X719 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X720 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X721 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X722 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X723 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X724 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X725 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X726 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X727 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X728 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X729 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X730 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X731 a_n11737_n14973# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X732 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X733 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X734 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X735 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X736 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X737 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X738 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X739 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X740 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X741 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X742 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X743 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X744 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X745 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X746 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X747 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X748 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X749 AVDD IREF a_n11737_n15980# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X750 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X751 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X752 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X753 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X754 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X755 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X756 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X757 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X758 AVSS a_n11737_n15980# a_n6139_n21443# AVSS nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X759 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X760 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X761 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X762 a_n13990_n5465# a_n11737_n15980# VOUT AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X763 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X764 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X765 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X766 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X767 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X768 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X769 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X770 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X771 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X772 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X773 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X774 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X775 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X776 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X777 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X778 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X779 AVDD IREF IREF AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X780 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X781 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X782 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X783 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X784 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X785 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X786 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X787 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X788 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X789 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X790 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X791 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X792 a_n11737_n14973# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X793 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X794 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X795 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X796 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X797 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X798 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X799 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X800 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X801 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X802 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X803 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X804 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X805 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X806 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X807 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X808 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X809 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X810 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X811 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X812 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X813 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X814 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X815 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X816 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X817 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X818 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X819 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X820 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X821 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X822 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X823 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X824 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X825 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X826 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X827 a_n11737_n14973# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X828 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X829 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X830 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X831 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X832 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X833 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X834 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X835 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X836 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X837 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X838 AVDD a_n11317_n20927# a_n1533_n17634# AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X839 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X840 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X841 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X842 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X843 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X844 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X845 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X846 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X847 a_5396_n6451# a_n11737_n15980# a_n13990_n6451# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X848 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X849 a_5396_n6451# a_n11737_n15980# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X850 a_n6139_n20267# a_n11737_n15980# a_n11737_n15980# AVSS nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X851 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X852 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X853 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X854 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X855 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X856 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X857 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X858 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X859 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X860 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X861 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X862 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X863 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X864 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X865 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X866 IREF IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X867 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X868 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X869 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X870 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X871 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X872 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X873 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X874 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X875 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X876 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X877 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X878 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X879 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X880 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X881 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X882 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X883 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X884 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X885 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X886 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X887 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X888 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X889 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X890 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X891 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X892 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X893 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X894 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X895 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X896 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X897 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X898 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X899 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X900 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X901 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X902 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X903 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X904 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X905 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X906 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X907 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X908 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X909 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X910 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X911 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X912 AVDD IREF a_n11737_n14973# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X913 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X914 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X915 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X916 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X917 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X918 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X919 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X920 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X921 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X922 a_n5579_n20820# a_n11737_n15980# a_n6139_n20820# AVSS nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X923 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X924 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X925 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X926 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X927 a_n13990_n5465# a_n11737_n15980# VOUT AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X928 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X929 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X930 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X931 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X932 a_n13990_n5465# a_n11737_n15980# VOUT AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X933 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X934 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X935 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X936 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X937 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X938 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X939 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X940 a_n11317_n20927# a_n11317_n20927# a_n965_n15598# AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.78p ps=3.7u w=1.2u l=2u
X941 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X942 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X943 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X944 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X945 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X946 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X947 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X948 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X949 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X950 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X951 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X952 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X953 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X954 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X955 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X956 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X957 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X958 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X959 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X960 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X961 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X962 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X963 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X964 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X965 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X966 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X967 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X968 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X969 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X970 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X971 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X972 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X973 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X974 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X975 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X976 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X977 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X978 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X979 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X980 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X981 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X982 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X983 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X984 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X985 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X986 a_n11737_n14973# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X987 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X988 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X989 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X990 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X991 AVDD IREF IREF AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X992 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X993 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X994 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X995 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X996 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X997 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X998 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X999 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1000 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1001 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1002 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1003 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1004 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1005 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1006 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1007 a_n11737_n15980# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1008 AVDD IREF IREF AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1009 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1010 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1011 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1012 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1013 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1014 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1015 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1016 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1017 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1018 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1019 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1020 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1021 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1022 a_n13990_n6451# a_n11737_n15980# a_5396_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1023 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1024 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1025 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1026 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1027 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1028 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1029 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1030 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1031 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1032 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1033 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1034 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1035 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1036 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1037 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1038 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1039 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1040 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1041 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1042 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1043 AVDD IREF a_n11737_n15980# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1044 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1045 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1046 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1047 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1048 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1049 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1050 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1051 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1052 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1053 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1054 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1055 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1056 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1057 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1058 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1059 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1060 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1061 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1062 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1063 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1064 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1065 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1066 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1067 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1068 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1069 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1070 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1071 a_n11737_n14973# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1072 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1073 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1074 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1075 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1076 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1077 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1078 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1079 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1080 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1081 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1082 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1083 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1084 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1085 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1086 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1087 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1088 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1089 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1090 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1091 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1092 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1093 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1094 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1095 AVSS a_n11737_n14973# a_n11317_n20927# AVSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X1096 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1097 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1098 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1099 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1100 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1101 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1102 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1103 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1104 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1105 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1106 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1107 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1108 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1109 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1110 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1111 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1112 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1113 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1114 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1115 VOUT a_n11737_n15980# a_n13990_n5465# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1116 VOUT a_n11737_n15980# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1117 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1118 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1119 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1120 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1121 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1122 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1123 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1124 AVSS a_n11737_n14973# a_n11737_n14973# AVSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X1125 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1126 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1127 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1128 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1129 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1130 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1131 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1132 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1133 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1134 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1135 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1136 a_n11737_n15980# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1137 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1138 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1139 AVDD IREF a_n11737_n14973# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1140 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1141 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1142 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1143 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1144 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1145 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1146 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1147 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1148 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1149 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1150 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1151 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1152 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1153 VOUT a_n11737_n15980# a_n13990_n5465# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1154 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1155 AVDD IREF a_n11737_n14973# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1156 VOUT a_n11737_n15980# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1157 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1158 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1159 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1160 AVDD IREF a_n11737_n15980# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1161 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1162 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1163 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1164 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1165 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1166 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1167 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1168 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1169 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X1170 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1171 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1172 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1173 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1174 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1175 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1176 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X1177 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1178 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1179 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1180 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1181 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1182 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1183 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1184 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1185 a_n13990_n6451# a_n11737_n15980# a_5396_n6451# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1186 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1187 a_n13990_n6451# a_n11737_n15980# a_5396_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1188 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1189 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1190 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1191 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1192 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1193 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1194 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1195 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1196 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1197 a_n11737_n15980# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1198 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1199 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1200 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1201 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1202 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1203 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1204 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1205 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1206 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1207 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1208 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1209 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1210 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1211 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1212 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1213 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1214 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1215 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1216 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1217 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1218 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1219 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1220 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1221 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1222 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X1223 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1224 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1225 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1226 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1227 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X1228 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1229 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1230 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1231 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1232 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1233 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1234 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1235 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1236 VOUT a_n11737_n15980# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1237 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1238 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1239 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1240 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1241 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1242 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1243 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1244 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1245 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1246 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1247 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1248 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1249 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1250 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1251 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1252 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1253 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1254 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1255 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1256 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1257 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1258 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1259 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1260 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1261 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1262 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1263 IREF IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1264 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1265 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1266 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1267 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1268 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1269 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1270 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1271 IREF IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1272 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1273 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1274 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1275 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1276 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1277 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1278 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1279 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1280 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1281 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1282 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1283 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1284 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1285 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1286 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1287 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1288 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1289 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1290 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1291 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1292 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1293 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1294 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1295 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1296 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1297 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1298 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1299 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1300 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1301 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1302 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1303 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1304 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1305 a_n13990_n6451# a_n11737_n15980# a_5396_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1306 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1307 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1308 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1309 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1310 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1311 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1312 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1313 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1314 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1315 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1316 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1317 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1318 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1319 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1320 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1321 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1322 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1323 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1324 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1325 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1326 a_n11737_n15980# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1327 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1328 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1329 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1330 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1331 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1332 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1333 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1334 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1335 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1336 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1337 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1338 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1339 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1340 AVDD IREF IREF AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1341 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1342 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1343 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1344 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1345 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1346 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1347 AVDD IREF IREF AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1348 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1349 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1350 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1351 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X1352 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1353 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1354 a_n13990_n6451# a_n11737_n15980# a_5396_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1355 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1356 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1357 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1358 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1359 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1360 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1361 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1362 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1363 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1364 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1365 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1366 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1367 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1368 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1369 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1370 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1371 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1372 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1373 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1374 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1375 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1376 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1377 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1378 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1379 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1380 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1381 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1382 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1383 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1384 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1385 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1386 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1387 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1388 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1389 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1390 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1391 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1392 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1393 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1394 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1395 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1396 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1397 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1398 AVDD IREF a_n11737_n15980# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1399 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1400 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1401 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1402 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1403 a_5396_n6451# a_n11737_n15980# a_n13990_n6451# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1404 a_5396_n6451# a_n11737_n15980# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1405 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1406 AVSS a_n11737_n14973# a_n13990_n6451# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1407 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1408 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1409 AVDD IREF a_n11737_n15980# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1410 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1411 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1412 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1413 a_n5579_n20820# a_n11737_n15980# a_n6139_n20267# AVSS nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X1414 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1415 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1416 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1417 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1418 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1419 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1420 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1421 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1422 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1423 a_n1533_n16909# a_n11317_n20927# a_n2101_n16909# AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X1424 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1425 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1426 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1427 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1428 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1429 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1430 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1431 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1432 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1433 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1434 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1435 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1436 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1437 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1438 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1439 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1440 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1441 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1442 VOUT a_n11737_n15980# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1443 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1444 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1445 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1446 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1447 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1448 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1449 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1450 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1451 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1452 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1453 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1454 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1455 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1456 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1457 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1458 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1459 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1460 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1461 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1462 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1463 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1464 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1465 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1466 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1467 AVDD IREF a_n11737_n15980# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1468 a_n11317_n20927# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X1469 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1470 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1471 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1472 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1473 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1474 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1475 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1476 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1477 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1478 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1479 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1480 AVDD IREF a_n11737_n14973# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1481 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1482 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1483 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1484 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1485 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1486 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1487 IREF IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1488 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1489 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1490 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1491 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1492 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1493 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1494 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1495 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1496 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1497 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1498 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1499 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1500 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1501 AVSS a_n11737_n14973# a_n13990_n5465# AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1502 a_n2101_n16909# a_n11317_n20927# a_n2631_n17634# AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X1503 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1504 a_5396_9163# a_n11317_n20927# VOUT AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1505 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1506 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1507 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1508 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1509 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1510 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1511 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1512 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1513 a_n13990_8177# VP a_n13990_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1514 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1515 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1516 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1517 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1518 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1519 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1520 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1521 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1522 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1523 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1524 AVDD IREF IREF AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1525 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1526 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1527 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1528 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1529 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1530 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1531 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1532 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1533 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1534 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1535 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1536 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1537 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1538 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1539 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1540 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1541 a_n11737_n15980# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1542 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1543 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1544 a_n11737_n14973# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1545 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1546 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1547 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1548 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1549 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1550 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1551 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1552 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1553 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1554 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1555 a_n11737_n14973# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1556 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1557 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1558 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1559 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1560 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1561 AVDD IREF IREF AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1562 a_n13990_n6451# VP a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1563 a_n13990_n6451# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1564 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1565 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X1566 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1567 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1568 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1569 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1570 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1571 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1572 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1573 a_n13990_8177# VN a_n13990_n5465# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1574 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1575 AVDD a_5396_n6451# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1576 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1577 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1578 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1579 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1580 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1581 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1582 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1583 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1584 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1585 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1586 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1587 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1588 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1589 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1590 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1591 AVSS AVSS AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1592 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1593 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1594 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1595 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1596 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1597 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1598 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1599 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1600 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1601 a_5396_8177# a_n11317_n20927# a_5396_n6451# AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1602 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1603 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1604 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1605 AVDD IREF a_n13990_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1606 a_n11737_n14973# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1607 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1608 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1609 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1610 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1611 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1612 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1613 VOUT a_n11317_n20927# a_5396_9163# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1614 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1615 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1616 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1617 AVSS AVSS AVSS AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1618 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1619 AVDD AVDD AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1620 a_n13990_n5465# VN a_n13990_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1621 a_5396_9163# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1622 a_n13990_n5465# a_n11737_n14973# AVSS AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1623 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1624 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1625 AVDD a_5396_n6451# a_5396_8177# AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1626 a_n13990_8177# IREF AVDD AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1627 AVDD AVDD AVDD AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1628 a_5396_n6451# a_n11317_n20927# a_5396_8177# AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1629 a_5396_8177# a_5396_n6451# AVDD AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
.ends

