** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/DiffP_pfets.sch
.subckt DiffP_pfets D1 D2 G1 G2 S B
*.PININFO D1:B D2:B G1:B G2:B S:B B:B
M1 net4 G1 S B pfet_03v3 L=2u W=2u nf=1 m=1
M2 net5 G2 S B pfet_03v3 L=2u W=2u nf=1 m=1
M5 net3 G1 S B pfet_03v3 L=2u W=2u nf=1 m=1
M6 net2 G1 S B pfet_03v3 L=2u W=2u nf=1 m=1
M7 net1 G1 S B pfet_03v3 L=2u W=2u nf=1 m=1
M8 D1 G1 net4 B pfet_03v3 L=2u W=2u nf=1 m=1
M9 D1 G1 net3 B pfet_03v3 L=2u W=2u nf=1 m=1
M10 D1 G1 net2 B pfet_03v3 L=2u W=2u nf=1 m=1
M11 D1 G1 net1 B pfet_03v3 L=2u W=2u nf=1 m=1
M12 net6 G2 S B pfet_03v3 L=2u W=2u nf=1 m=1
M15 D2 G2 net5 B pfet_03v3 L=2u W=2u nf=1 m=1
M16 D2 G2 net6 B pfet_03v3 L=2u W=2u nf=1 m=1
M19 net7 G2 S B pfet_03v3 L=2u W=2u nf=1 m=1
M20 net8 G2 S B pfet_03v3 L=2u W=2u nf=1 m=1
M21 D2 G2 net7 B pfet_03v3 L=2u W=2u nf=1 m=1
M22 D2 G2 net8 B pfet_03v3 L=2u W=2u nf=1 m=1
M3[1] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[2] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[3] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[4] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[5] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[6] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[7] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[8] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[9] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[10] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[11] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[12] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[13] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[14] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[15] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[16] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[17] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[18] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[19] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[20] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[21] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[22] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[23] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[24] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[25] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[26] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[27] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[28] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[29] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[30] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[31] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[32] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
.ends
.end
