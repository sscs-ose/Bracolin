* Extracted by KLayout with GF180MCU LVS runset on : 04/01/2024 22:27

.SUBCKT Filter_TOP A2 B2 AVDD|AVSS|VDD|VSS B1|VOUT CMOUTP CMOUTN ISBCS ISBCS2
+ IREF VP A1|VN gf180mcu_gnd
M$1 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$4 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$5 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$6 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$7 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$8 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$9 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$10 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$11 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$12 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$13 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$14 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$15 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$16 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$17 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$18 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$19 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$20 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$21 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$22 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$23 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$24 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$25 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$26 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$27 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$28 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$29 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$30 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$31 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$32 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$33 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$34 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$35 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$36 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$37 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$38 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$39 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$40 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$41 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$42 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$43 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$44 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$45 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$46 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$47 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$48 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$49 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$50 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$51 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$52 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$53 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$54 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$55 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$56 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$57 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$58 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$59 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$60 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$61 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$62 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$63 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$64 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$65 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$66 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$67 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$68 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$69 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$70 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$71 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$72 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$73 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$74 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$75 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$76 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$77 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$78 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$79 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$80 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$81 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$82 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$83 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$84 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$85 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$86 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$87 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$88 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$89 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$90 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$91 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$92 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$93 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$94 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$95 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$96 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$97 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$98 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$99 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$100 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$101 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$102 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$103 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$104 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$105 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$106 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$107 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$108 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$109 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$110 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$111 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$112 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$113 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$114 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$115 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$116 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$117 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$118 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$119 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$120 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$121 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$122 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$123 \$135 \$172 \$917 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$124 AVDD|AVSS|VDD|VSS \$172 \$135 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$125 \$136 \$172 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$126 \$172 \$172 \$136 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$127 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$128 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$129 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$130 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$131 \$137 \$24 \$1 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$132 \$138 \$24 \$137 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$133 \$139 \$24 \$115 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$134 A2 \$24 \$139 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$135 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$136 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$137 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$138 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$139 \$141 \$173 \$24 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$140 \$29 \$173 \$141 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$141 \$142 \$258 \$29 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$142 \$257 \$258 \$142 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$143 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$144 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$145 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$146 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$147 \$143 \$174 \$919 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$148 AVDD|AVSS|VDD|VSS \$174 \$143 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$149 \$144 \$174 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$150 \$174 \$174 \$144 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$151 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$152 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$153 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$154 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$155 \$145 \$25 \$2 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$156 \$146 \$25 \$145 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$157 \$147 \$25 \$116 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$158 \$1 \$25 \$147 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$159 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$160 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$161 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$162 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$163 \$148 \$175 \$25 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$164 \$30 \$175 \$148 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$165 \$149 \$260 \$30 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$166 \$259 \$260 \$149 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$167 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$168 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$169 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$170 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$171 \$150 \$176 \$921 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$172 AVDD|AVSS|VDD|VSS \$176 \$150 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$173 \$151 \$176 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$174 \$176 \$176 \$151 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$175 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$176 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$177 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$178 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$179 \$152 \$26 \$3 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$180 \$153 \$26 \$152 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$181 \$154 \$26 \$117 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$182 \$2 \$26 \$154 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$183 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$184 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$185 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$186 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$187 \$155 \$177 \$26 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$188 \$31 \$177 \$155 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$189 \$156 \$262 \$31 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$190 \$261 \$262 \$156 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$191 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$192 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$193 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$194 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$195 \$157 \$178 \$923 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$196 AVDD|AVSS|VDD|VSS \$178 \$157 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$197 \$158 \$178 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$198 \$178 \$178 \$158 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$199 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$200 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$201 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$202 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$203 \$159 \$27 \$4 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$204 \$160 \$27 \$159 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$205 \$161 \$27 \$118 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$206 \$3 \$27 \$161 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$207 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$208 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$209 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$210 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$211 \$162 \$179 \$27 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$212 \$32 \$179 \$162 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$213 \$163 \$264 \$32 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$214 \$263 \$264 \$163 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$215 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$216 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$217 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$218 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$219 \$164 \$180 \$925 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$220 AVDD|AVSS|VDD|VSS \$180 \$164 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$221 \$165 \$180 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$222 \$180 \$180 \$165 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$223 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$224 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$225 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$226 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$227 \$167 \$28 B2 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$228 \$168 \$28 \$167 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$229 \$169 \$28 \$119 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$230 \$4 \$28 \$169 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$231 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$232 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$233 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$234 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$235 \$170 \$181 \$28 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$236 \$33 \$181 \$170 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$237 \$171 \$266 \$33 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$238 \$265 \$266 \$171 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$239 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$240 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$241 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$242 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$243 \$307 \$172 \$172 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$244 AVDD|AVSS|VDD|VSS \$172 \$307 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$245 \$308 \$172 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$246 \$917 \$172 \$308 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$247 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$248 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$249 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$250 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$251 \$309 \$24 \$173 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$252 AVDD|AVSS|VDD|VSS \$24 \$309 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$253 \$310 \$24 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$254 \$173 \$24 \$310 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$255 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$256 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$257 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$258 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$259 \$311 \$258 \$257 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$260 \$29 \$258 \$311 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$261 \$312 \$173 \$29 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$262 \$24 \$173 \$312 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$263 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$264 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$265 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$266 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$267 \$313 \$174 \$174 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$268 AVDD|AVSS|VDD|VSS \$174 \$313 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$269 \$314 \$174 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$270 \$919 \$174 \$314 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$271 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$272 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$273 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$274 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$275 \$315 \$25 \$175 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$276 AVDD|AVSS|VDD|VSS \$25 \$315 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$277 \$316 \$25 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$278 \$175 \$25 \$316 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$279 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$280 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$281 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$282 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$283 \$317 \$260 \$259 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$284 \$30 \$260 \$317 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$285 \$318 \$175 \$30 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$286 \$25 \$175 \$318 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$287 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$288 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$289 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$290 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$291 \$319 \$176 \$176 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$292 AVDD|AVSS|VDD|VSS \$176 \$319 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$293 \$320 \$176 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$294 \$921 \$176 \$320 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$295 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$296 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$297 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$298 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$299 \$321 \$26 \$177 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$300 AVDD|AVSS|VDD|VSS \$26 \$321 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$301 \$322 \$26 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$302 \$177 \$26 \$322 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$303 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$304 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$305 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$306 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$307 \$323 \$262 \$261 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$308 \$31 \$262 \$323 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$309 \$324 \$177 \$31 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$310 \$26 \$177 \$324 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$311 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$312 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$313 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$314 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$315 \$325 \$178 \$178 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$316 AVDD|AVSS|VDD|VSS \$178 \$325 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$317 \$326 \$178 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$318 \$923 \$178 \$326 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$319 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$320 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$321 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$322 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$323 \$327 \$27 \$179 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$324 AVDD|AVSS|VDD|VSS \$27 \$327 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$325 \$328 \$27 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$326 \$179 \$27 \$328 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$327 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$328 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$329 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$330 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$331 \$329 \$264 \$263 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$332 \$32 \$264 \$329 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$333 \$330 \$179 \$32 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$334 \$27 \$179 \$330 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$335 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$336 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$337 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$338 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$339 \$331 \$180 \$180 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$340 AVDD|AVSS|VDD|VSS \$180 \$331 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$341 \$332 \$180 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$342 \$925 \$180 \$332 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$343 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$344 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$345 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$346 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$347 \$333 \$28 \$181 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$348 AVDD|AVSS|VDD|VSS \$28 \$333 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$349 \$334 \$28 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$350 \$181 \$28 \$334 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$351 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$352 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$353 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$354 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$355 \$335 \$266 \$265 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$356 \$33 \$266 \$335 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$357 \$336 \$181 \$33 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$358 \$28 \$181 \$336 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$359 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$360 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$361 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$362 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$363 \$442 \$172 \$917 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$364 AVDD|AVSS|VDD|VSS \$172 \$442 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$365 \$443 \$172 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$366 \$172 \$172 \$443 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$367 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$368 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$369 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$370 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$371 \$444 \$24 \$173 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$372 AVDD|AVSS|VDD|VSS \$24 \$444 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$373 \$445 \$24 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$374 \$173 \$24 \$445 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$375 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$376 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$377 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$378 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$379 \$446 \$173 \$24 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$380 \$29 \$173 \$446 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$381 \$447 \$258 \$29 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$382 \$257 \$258 \$447 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$383 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$384 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$385 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$386 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$387 \$448 \$174 \$919 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$388 AVDD|AVSS|VDD|VSS \$174 \$448 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$389 \$449 \$174 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$390 \$174 \$174 \$449 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$391 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$392 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$393 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$394 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$395 \$450 \$25 \$175 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$396 AVDD|AVSS|VDD|VSS \$25 \$450 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$397 \$451 \$25 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$398 \$175 \$25 \$451 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$399 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$400 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$401 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$402 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$403 \$452 \$175 \$25 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$404 \$30 \$175 \$452 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$405 \$453 \$260 \$30 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$406 \$259 \$260 \$453 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$407 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$408 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$409 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$410 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$411 \$454 \$176 \$921 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$412 AVDD|AVSS|VDD|VSS \$176 \$454 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$413 \$455 \$176 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$414 \$176 \$176 \$455 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$415 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$416 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$417 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$418 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$419 \$456 \$26 \$177 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$420 AVDD|AVSS|VDD|VSS \$26 \$456 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$421 \$457 \$26 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$422 \$177 \$26 \$457 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$423 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$424 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$425 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$426 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$427 \$458 \$177 \$26 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$428 \$31 \$177 \$458 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$429 \$459 \$262 \$31 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$430 \$261 \$262 \$459 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$431 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$432 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$433 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$434 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$435 \$460 \$178 \$923 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$436 AVDD|AVSS|VDD|VSS \$178 \$460 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$437 \$461 \$178 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$438 \$178 \$178 \$461 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$439 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$440 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$441 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$442 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$443 \$462 \$27 \$179 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$444 AVDD|AVSS|VDD|VSS \$27 \$462 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$445 \$463 \$27 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$446 \$179 \$27 \$463 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$447 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$448 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$449 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$450 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$451 \$464 \$179 \$27 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$452 \$32 \$179 \$464 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$453 \$465 \$264 \$32 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$454 \$263 \$264 \$465 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$455 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$456 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$457 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$458 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$459 \$466 \$180 \$925 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$460 AVDD|AVSS|VDD|VSS \$180 \$466 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$461 \$467 \$180 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$462 \$180 \$180 \$467 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$463 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$464 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$465 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$466 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$467 \$468 \$28 \$181 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$468 AVDD|AVSS|VDD|VSS \$28 \$468 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$469 \$469 \$28 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$470 \$181 \$28 \$469 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$471 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$472 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$473 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$474 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$475 \$470 \$181 \$28 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$476 \$33 \$181 \$470 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$477 \$471 \$266 \$33 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$478 \$265 \$266 \$471 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$479 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$480 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$481 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$482 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$483 \$587 \$172 \$172 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$484 AVDD|AVSS|VDD|VSS \$172 \$587 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$485 \$588 \$172 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$486 \$917 \$172 \$588 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$487 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$488 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$489 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$490 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$491 \$589 \$24 A2 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$492 \$115 \$24 \$589 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$493 \$590 \$24 \$138 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$494 \$1 \$24 \$590 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$495 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$496 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$497 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$498 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$499 \$591 \$258 \$257 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$500 \$29 \$258 \$591 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$501 \$592 \$173 \$29 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$502 \$24 \$173 \$592 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$503 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$504 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$505 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$506 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$507 \$593 \$174 \$174 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$508 AVDD|AVSS|VDD|VSS \$174 \$593 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$509 \$594 \$174 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$510 \$919 \$174 \$594 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$511 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$512 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$513 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$514 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$515 \$595 \$25 \$1 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$516 \$116 \$25 \$595 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$517 \$596 \$25 \$146 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$518 \$2 \$25 \$596 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$519 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$520 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$521 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$522 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$523 \$597 \$260 \$259 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$524 \$30 \$260 \$597 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$525 \$598 \$175 \$30 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$526 \$25 \$175 \$598 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$527 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$528 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$529 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$530 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$531 \$599 \$176 \$176 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$532 AVDD|AVSS|VDD|VSS \$176 \$599 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$533 \$600 \$176 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$534 \$921 \$176 \$600 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$535 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$536 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$537 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$538 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$539 \$601 \$26 \$2 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$540 \$117 \$26 \$601 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$541 \$602 \$26 \$153 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$542 \$3 \$26 \$602 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$543 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$544 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$545 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$546 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$547 \$603 \$262 \$261 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$548 \$31 \$262 \$603 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$549 \$604 \$177 \$31 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$550 \$26 \$177 \$604 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$551 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$552 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$553 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$554 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$555 \$605 \$178 \$178 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$556 AVDD|AVSS|VDD|VSS \$178 \$605 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$557 \$606 \$178 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$558 \$923 \$178 \$606 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$559 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$560 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$561 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$562 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$563 \$607 \$27 \$3 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$564 \$118 \$27 \$607 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$565 \$608 \$27 \$160 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$566 \$4 \$27 \$608 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$567 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$568 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$569 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$570 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$571 \$609 \$264 \$263 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$572 \$32 \$264 \$609 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$573 \$610 \$179 \$32 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$574 \$27 \$179 \$610 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$575 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$576 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$577 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$578 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$579 \$611 \$180 \$180 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$580 AVDD|AVSS|VDD|VSS \$180 \$611 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$581 \$612 \$180 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$582 \$925 \$180 \$612 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$583 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$584 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$585 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$586 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$587 \$613 \$28 \$4 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$588 \$119 \$28 \$613 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$589 \$614 \$28 \$168 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$590 B2 \$28 \$614 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$591 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$592 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$593 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$594 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$595 \$615 \$266 \$265 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$596 \$33 \$266 \$615 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$597 \$616 \$181 \$33 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$598 \$28 \$181 \$616 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$599 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$600 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$601 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$602 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$603 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$604 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$605 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$606 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$607 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$608 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$609 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$610 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$611 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$612 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$613 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$614 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$615 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$616 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$617 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$618 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$619 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$620 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$621 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$622 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$623 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$624 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$625 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$626 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$627 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$628 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$629 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$630 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$631 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$632 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$633 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$634 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$635 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$636 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$637 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$638 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$639 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$640 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$641 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$642 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$643 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$644 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$645 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$646 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$647 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$648 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$649 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$650 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$651 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$652 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$653 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$654 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$655 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$656 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$657 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$658 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$659 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$660 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$661 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$662 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$663 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$664 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$665 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$666 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$667 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$668 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$669 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$670 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$671 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$672 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$673 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$674 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$675 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$676 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$677 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$678 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$679 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$680 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$681 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$682 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$683 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$684 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$685 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$686 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$687 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$688 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$689 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$690 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$691 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$692 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$693 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$694 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$695 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$696 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$697 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$698 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$699 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$700 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$701 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$702 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$703 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$704 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$705 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$706 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$707 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$708 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$709 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$710 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$711 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$712 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$713 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$714 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$715 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$716 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$717 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$718 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$719 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$720 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$721 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$722 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$723 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$724 \$1584 \$1573 \$1583 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$725 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$726 \$1671 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$727 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$728 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$729 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$730 \$1585 \$1573 \$1584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$731 \$1586 \$1573 \$1585 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$732 \$1587 \$1573 \$1586 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$733 \$1672 \$1573 \$1671 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$734 \$1673 \$1573 \$1672 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$735 \$1674 \$1573 \$1673 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$736 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$737 AVDD|AVSS|VDD|VSS \$1573 \$1587 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$738 \$1675 \$1573 \$1674 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$739 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$740 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$741 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$742 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$743 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$744 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$745 \$1676 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$746 \$1589 \$1573 \$1588 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$747 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$748 \$1590 \$1573 \$1589 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$749 \$1591 \$1573 \$1590 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$750 \$1592 \$1573 \$1591 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$751 \$1677 \$1573 \$1676 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$752 \$1678 \$1573 \$1677 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$753 \$1679 \$1573 \$1678 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$754 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$755 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$756 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$757 AVDD|AVSS|VDD|VSS \$1573 \$1592 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$758 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$759 \$1680 \$1573 \$1679 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$760 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$761 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$762 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$763 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$764 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$765 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$766 \$1681 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$767 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$768 \$1594 \$1573 \$1593 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$769 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$770 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$771 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$772 \$1595 \$1573 \$1594 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$773 \$1596 \$1573 \$1595 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$774 \$1597 \$1573 \$1596 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$775 \$1682 \$1573 \$1681 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$776 \$1683 \$1573 \$1682 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$777 \$1684 \$1573 \$1683 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$778 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$779 AVDD|AVSS|VDD|VSS \$1573 \$1597 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$780 \$1685 \$1573 \$1684 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$781 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$782 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$783 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$784 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$785 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$786 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$787 \$1686 \$1574 \$173 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P
+ PS=5.3U PD=5.3U
M$788 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$789 \$1599 \$1574 \$1598 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$790 \$1687 \$1574 \$1686 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$791 \$1688 \$1574 \$1687 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$792 \$1689 \$1574 \$1688 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$793 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$794 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$795 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$796 \$1600 \$1574 \$1599 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$797 \$1601 \$1574 \$1600 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$798 \$1602 \$1574 \$1601 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$799 \$1603 \$1574 \$1602 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$800 \$1690 \$1574 \$1689 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$801 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$802 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$803 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$804 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$805 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$806 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$807 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$808 \$1691 \$1574 \$175 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P
+ PS=5.3U PD=5.3U
M$809 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$810 \$1605 \$1574 \$1604 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$811 \$1606 \$1574 \$1605 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$812 \$1607 \$1574 \$1606 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$813 \$1608 \$1574 \$1607 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$814 \$1692 \$1574 \$1691 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$815 \$1693 \$1574 \$1692 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$816 \$1694 \$1574 \$1693 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$817 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$818 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$819 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$820 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$821 \$1609 \$1574 \$1608 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$822 \$1695 \$1574 \$1694 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$823 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$824 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$825 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$826 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$827 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$828 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$829 \$1611 \$1574 \$1610 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$830 \$1696 \$1574 \$177 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P
+ PS=5.3U PD=5.3U
M$831 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$832 \$1697 \$1574 \$1696 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$833 \$1698 \$1574 \$1697 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$834 \$1699 \$1574 \$1698 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$835 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$836 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$837 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$838 \$1612 \$1574 \$1611 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$839 \$1613 \$1574 \$1612 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$840 \$1614 \$1574 \$1613 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$841 \$1700 \$1574 \$1699 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$842 \$1615 \$1574 \$1614 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$843 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$844 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$845 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$846 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$847 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$848 \$1821 \$1573 \$1820 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$849 \$1822 \$1573 \$1821 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$850 \$1823 \$1573 \$1822 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$851 \$1824 \$1573 \$1823 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$852 \$1675 \$1573 \$1824 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$853 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$854 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$855 \$1826 \$1573 \$1825 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$856 \$1827 \$1573 \$1826 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$857 \$1828 \$1573 \$1827 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$858 \$1829 \$1573 \$1828 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$859 \$1680 \$1573 \$1829 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$860 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$861 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$862 \$1831 \$1573 \$1830 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$863 \$1832 \$1573 \$1831 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$864 \$1833 \$1573 \$1832 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$865 \$1834 \$1573 \$1833 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$866 \$1685 \$1573 \$1834 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$867 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$868 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$869 \$1836 \$1574 \$1835 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$870 \$1837 \$1574 \$1836 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$871 \$1838 \$1574 \$1837 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$872 \$1839 \$1574 \$1838 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$873 \$1690 \$1574 \$1839 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$874 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$875 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$876 \$1841 \$1574 \$1840 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$877 \$1842 \$1574 \$1841 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$878 \$1843 \$1574 \$1842 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$879 \$1844 \$1574 \$1843 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$880 \$1695 \$1574 \$1844 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$881 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$882 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$883 \$1846 \$1574 \$1845 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$884 \$1847 \$1574 \$1846 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$885 \$1848 \$1574 \$1847 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$886 \$1849 \$1574 \$1848 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$887 \$1700 \$1574 \$1849 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$888 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$889 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$890 \$1976 \$1573 \$1820 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$891 \$1977 \$1573 \$1976 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$892 \$1978 \$1573 \$1977 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$893 \$1979 \$1573 \$1978 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$894 \$1980 \$1573 \$1979 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$895 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$896 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$897 \$1981 \$1573 \$1825 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$898 \$1982 \$1573 \$1981 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$899 \$1983 \$1573 \$1982 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$900 \$1984 \$1573 \$1983 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$901 \$1985 \$1573 \$1984 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$902 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$903 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$904 \$1986 \$1573 \$1830 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$905 \$1987 \$1573 \$1986 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$906 \$1988 \$1573 \$1987 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$907 \$1989 \$1573 \$1988 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$908 \$1990 \$1573 \$1989 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$909 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$910 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$911 \$1991 \$1574 \$1835 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$912 \$1992 \$1574 \$1991 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$913 \$1993 \$1574 \$1992 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$914 \$1994 \$1574 \$1993 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$915 \$1995 \$1574 \$1994 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$916 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$917 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$918 \$1996 \$1574 \$1840 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$919 \$1997 \$1574 \$1996 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$920 \$1998 \$1574 \$1997 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$921 \$1999 \$1574 \$1998 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$922 \$2000 \$1574 \$1999 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$923 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$924 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$925 \$2001 \$1574 \$1845 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$926 \$2002 \$1574 \$2001 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$927 \$2003 \$1574 \$2002 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$928 \$2004 \$1574 \$2003 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$929 \$2005 \$1574 \$2004 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$930 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$931 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$932 \$2147 \$1573 \$1583 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$933 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$934 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$935 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$936 \$2149 \$1573 \$2148 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$937 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$938 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$939 \$2150 \$1573 \$1588 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$940 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$941 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$942 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$943 \$2152 \$1573 \$2151 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$944 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$945 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$946 \$2153 \$1573 \$1593 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$947 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$948 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$949 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$950 \$2154 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$951 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$952 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$953 \$2155 \$1574 \$1598 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$954 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$955 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$956 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$957 \$2156 \$1574 \$1603 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$958 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$959 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$960 \$2157 \$1574 \$1604 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$961 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$962 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$963 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$964 \$2158 \$1574 \$1609 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$965 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$966 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$967 \$2159 \$1574 \$1610 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$968 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$969 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$970 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$971 \$2160 \$1574 \$1615 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$972 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$973 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$974 \$2147 \$1573 \$2290 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$975 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$976 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$977 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$978 \$2149 \$1573 \$2291 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$979 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$980 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$981 \$2150 \$1573 \$2292 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$982 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$983 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$984 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$985 \$2152 \$1573 \$2293 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$986 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$987 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$988 \$2153 \$1573 \$2294 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$989 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$990 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$991 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$992 \$2154 \$1573 \$2295 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$993 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$994 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$995 \$2155 \$1574 \$2296 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$996 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$997 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$998 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$999 \$2156 \$1574 \$29 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P
+ PS=5.3U PD=5.3U
M$1000 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1001 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1002 \$2157 \$1574 \$2297 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1003 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1004 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1005 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1006 \$2158 \$1574 \$30 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P
+ PS=5.3U PD=5.3U
M$1007 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1008 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1009 \$2159 \$1574 \$2298 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1010 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1011 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1012 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1013 \$2160 \$1574 \$31 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P
+ PS=5.3U PD=5.3U
M$1014 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1015 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1016 \$2447 \$1573 \$2446 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1017 \$2448 \$1573 \$2447 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1018 \$2449 \$1573 \$2448 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1019 \$2450 \$1573 \$2449 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1020 \$1980 \$1573 \$2450 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1021 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1022 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1023 \$2452 \$1573 \$2451 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1024 \$2453 \$1573 \$2452 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1025 \$2454 \$1573 \$2453 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1026 \$2455 \$1573 \$2454 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1027 \$1985 \$1573 \$2455 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1028 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1029 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1030 \$2457 \$1573 \$2456 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1031 \$2458 \$1573 \$2457 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1032 \$2459 \$1573 \$2458 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1033 \$2460 \$1573 \$2459 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1034 \$1990 \$1573 \$2460 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1035 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1036 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1037 \$2462 \$1574 \$2461 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1038 \$2463 \$1574 \$2462 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1039 \$2464 \$1574 \$2463 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1040 \$2465 \$1574 \$2464 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1041 \$1995 \$1574 \$2465 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1042 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1043 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1044 \$2467 \$1574 \$2466 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1045 \$2468 \$1574 \$2467 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1046 \$2469 \$1574 \$2468 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1047 \$2470 \$1574 \$2469 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1048 \$2000 \$1574 \$2470 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1049 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1050 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1051 \$2472 \$1574 \$2471 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1052 \$2473 \$1574 \$2472 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1053 \$2474 \$1574 \$2473 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1054 \$2475 \$1574 \$2474 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1055 \$2005 \$1574 \$2475 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1056 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1057 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1058 \$2648 \$1573 \$2446 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1059 \$2649 \$1573 \$2648 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1060 \$2650 \$1573 \$2649 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1061 \$2651 \$1573 \$2650 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1062 \$2652 \$1573 \$2651 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1063 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1064 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1065 \$2653 \$1573 \$2451 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1066 \$2654 \$1573 \$2653 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1067 \$2655 \$1573 \$2654 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1068 \$2656 \$1573 \$2655 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1069 \$2657 \$1573 \$2656 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1070 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1071 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1072 \$2658 \$1573 \$2456 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1073 \$2659 \$1573 \$2658 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1074 \$2660 \$1573 \$2659 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1075 \$2661 \$1573 \$2660 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1076 \$2662 \$1573 \$2661 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1077 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1078 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1079 \$2663 \$1574 \$2461 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1080 \$2664 \$1574 \$2663 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1081 \$2665 \$1574 \$2664 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1082 \$2666 \$1574 \$2665 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1083 \$2667 \$1574 \$2666 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1084 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1085 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1086 \$2668 \$1574 \$2466 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1087 \$2669 \$1574 \$2668 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1088 \$2670 \$1574 \$2669 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1089 \$2671 \$1574 \$2670 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1090 \$2672 \$1574 \$2671 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1091 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1092 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1093 \$2673 \$1574 \$2471 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1094 \$2674 \$1574 \$2673 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1095 \$2675 \$1574 \$2674 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1096 \$2676 \$1574 \$2675 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1097 \$2677 \$1574 \$2676 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1098 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1099 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1100 \$2960 \$1573 \$6258 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1101 \$2961 \$1573 \$2960 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1102 \$2962 \$1573 \$2961 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1103 \$2963 \$1573 \$2962 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1104 \$2652 \$1573 \$2963 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1105 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1106 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1107 \$2964 \$1573 \$6259 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1108 \$2965 \$1573 \$2964 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1109 \$2966 \$1573 \$2965 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1110 \$2967 \$1573 \$2966 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1111 \$2657 \$1573 \$2967 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1112 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1113 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1114 \$2969 \$1573 CMOUTP AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1115 \$2970 \$1573 \$2969 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1116 \$2971 \$1573 \$2970 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1117 \$2972 \$1573 \$2971 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1118 \$2662 \$1573 \$2972 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1119 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1120 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1121 \$2973 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1122 \$2974 \$1574 \$2973 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1123 \$2975 \$1574 \$2974 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1124 \$2976 \$1574 \$2975 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1125 \$2667 \$1574 \$2976 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1126 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1127 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1128 \$2977 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1129 \$2978 \$1574 \$2977 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1130 \$2979 \$1574 \$2978 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1131 \$2980 \$1574 \$2979 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1132 \$2672 \$1574 \$2980 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1133 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1134 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1135 \$2981 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1136 \$2982 \$1574 \$2981 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1137 \$2983 \$1574 \$2982 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1138 \$2984 \$1574 \$2983 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1139 \$2677 \$1574 \$2984 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1140 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1141 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1142 \$3235 \$1573 \$2290 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1143 \$3236 \$1573 \$3235 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1144 \$3237 \$1573 \$3236 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1145 \$3238 \$1573 \$3237 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1146 \$2291 \$1573 \$3238 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1147 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1148 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1149 \$3239 \$1573 \$2292 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1150 \$3240 \$1573 \$3239 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1151 \$3241 \$1573 \$3240 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1152 \$3242 \$1573 \$3241 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1153 \$2293 \$1573 \$3242 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1154 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1155 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1156 \$3243 \$1573 \$2294 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1157 \$3244 \$1573 \$3243 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1158 \$3245 \$1573 \$3244 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1159 \$3246 \$1573 \$3245 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1160 \$2295 \$1573 \$3246 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1161 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1162 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1163 \$3247 \$1574 \$2296 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1164 \$3248 \$1574 \$3247 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1165 \$3249 \$1574 \$3248 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1166 \$3250 \$1574 \$3249 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1167 AVDD|AVSS|VDD|VSS \$1574 \$3250 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1168 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1169 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1170 \$3251 \$1574 \$2297 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1171 \$3252 \$1574 \$3251 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1172 \$3253 \$1574 \$3252 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1173 \$3254 \$1574 \$3253 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1174 AVDD|AVSS|VDD|VSS \$1574 \$3254 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1175 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1176 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1177 \$3255 \$1574 \$2298 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1178 \$3256 \$1574 \$3255 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1179 \$3257 \$1574 \$3256 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1180 \$3258 \$1574 \$3257 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1181 AVDD|AVSS|VDD|VSS \$1574 \$3258 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1182 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1183 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1184 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1185 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1186 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1187 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1188 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1189 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1190 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1191 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1192 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1193 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1194 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1195 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1196 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1197 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1198 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1199 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1200 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1201 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1202 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1203 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1204 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1205 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1206 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1207 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1208 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1209 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1210 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1211 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1212 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1213 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1214 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1215 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1216 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1217 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1218 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1219 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1220 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1221 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1222 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1223 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1224 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1225 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1226 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1227 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1228 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1229 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1230 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1231 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1232 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1233 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1234 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1235 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1236 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1237 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1238 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1239 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1240 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1241 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1242 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1243 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1244 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1245 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1246 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1247 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1248 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1249 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1250 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1251 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1252 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1253 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1254 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1255 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1256 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1257 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1258 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1259 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1260 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1261 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1263 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1264 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1265 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1266 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1267 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1268 \$3563 \$1573 \$3562 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1269 \$3564 \$1573 \$3563 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1270 \$3565 \$1573 \$3564 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1271 \$3566 \$1573 \$3565 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1272 AVDD|AVSS|VDD|VSS \$1573 \$3566 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1273 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1274 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1275 \$3568 \$1573 \$3567 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1276 \$3569 \$1573 \$3568 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1277 \$3570 \$1573 \$3569 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1278 \$3571 \$1573 \$3570 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1279 AVDD|AVSS|VDD|VSS \$1573 \$3571 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1280 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1281 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1282 \$3573 \$1573 \$3572 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1283 \$3574 \$1573 \$3573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1284 \$3575 \$1573 \$3574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1285 \$3576 \$1573 \$3575 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1286 AVDD|AVSS|VDD|VSS \$1573 \$3576 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1287 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1288 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1289 \$3578 \$1574 \$3577 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1290 \$3579 \$1574 \$3578 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1291 \$3580 \$1574 \$3579 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1292 \$3581 \$1574 \$3580 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1293 \$3582 \$1574 \$3581 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1294 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1295 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1296 \$3584 \$1574 \$3583 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1297 \$3585 \$1574 \$3584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1298 \$3586 \$1574 \$3585 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1299 \$3587 \$1574 \$3586 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1300 \$3588 \$1574 \$3587 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1301 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1302 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1303 \$3590 \$1574 \$3589 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1304 \$3591 \$1574 \$3590 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1305 \$3592 \$1574 \$3591 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1306 \$3593 \$1574 \$3592 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1307 \$3594 \$1574 \$3593 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1308 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1309 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1310 \$3743 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1311 \$3744 \$1573 \$3743 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1312 \$3745 \$1573 \$3744 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1313 \$3746 \$1573 \$3745 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1314 \$3747 \$1573 \$3746 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1315 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1316 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1317 \$3748 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1318 \$3749 \$1573 \$3748 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1319 \$3750 \$1573 \$3749 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1320 \$3751 \$1573 \$3750 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1321 \$3752 \$1573 \$3751 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1322 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1323 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1324 \$3753 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1325 \$3754 \$1573 \$3753 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1326 \$3755 \$1573 \$3754 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1327 \$3756 \$1573 \$3755 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1328 \$3757 \$1573 \$3756 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1329 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1330 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1331 \$3758 \$1574 \$179 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1332 \$3759 \$1574 \$3758 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1333 \$3760 \$1574 \$3759 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1334 \$3761 \$1574 \$3760 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1335 \$3762 \$1574 \$3761 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1336 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1337 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1338 \$3763 \$1574 \$181 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1339 \$3764 \$1574 \$3763 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1340 \$3765 \$1574 \$3764 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1341 \$3766 \$1574 \$3765 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1342 \$3767 \$1574 \$3766 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1343 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1344 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1345 \$3768 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1346 \$3769 \$1574 \$3768 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1347 \$3770 \$1574 \$3769 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1348 \$3771 \$1574 \$3770 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1349 \$3772 \$1574 \$3771 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1350 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1351 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1352 \$3903 \$1573 \$3902 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1353 \$3904 \$1573 \$3903 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1354 \$3905 \$1573 \$3904 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1355 \$3906 \$1573 \$3905 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1356 \$3747 \$1573 \$3906 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1357 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1358 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1359 \$3908 \$1573 \$3907 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1360 \$3909 \$1573 \$3908 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1361 \$3910 \$1573 \$3909 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1362 \$3911 \$1573 \$3910 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1363 \$3752 \$1573 \$3911 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1364 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1365 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1366 \$3913 \$1573 \$3912 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1367 \$3914 \$1573 \$3913 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1368 \$3915 \$1573 \$3914 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1369 \$3916 \$1573 \$3915 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1370 \$3757 \$1573 \$3916 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1371 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1372 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1373 \$3918 \$1574 \$3917 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1374 \$3919 \$1574 \$3918 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1375 \$3920 \$1574 \$3919 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1376 \$3921 \$1574 \$3920 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1377 \$3762 \$1574 \$3921 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1378 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1379 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1380 \$3923 \$1574 \$3922 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1381 \$3924 \$1574 \$3923 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1382 \$3925 \$1574 \$3924 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1383 \$3926 \$1574 \$3925 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1384 \$3767 \$1574 \$3926 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1385 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1386 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1387 \$3928 \$1574 \$3927 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1388 \$3929 \$1574 \$3928 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1389 \$3930 \$1574 \$3929 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1390 \$3931 \$1574 \$3930 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1391 \$3772 \$1574 \$3931 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1392 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1393 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1394 \$4058 \$1573 \$3902 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1395 \$4059 \$1573 \$4058 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1396 \$4060 \$1573 \$4059 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1397 \$4061 \$1573 \$4060 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1398 \$4062 \$1573 \$4061 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1399 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1400 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1401 \$4063 \$1573 \$3907 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1402 \$4064 \$1573 \$4063 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1403 \$4065 \$1573 \$4064 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1404 \$4066 \$1573 \$4065 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1405 \$4067 \$1573 \$4066 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1406 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1407 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1408 \$4068 \$1573 \$3912 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1409 \$4069 \$1573 \$4068 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1410 \$4070 \$1573 \$4069 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1411 \$4071 \$1573 \$4070 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1412 \$4072 \$1573 \$4071 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1413 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1414 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1415 \$4073 \$1574 \$3917 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1416 \$4074 \$1574 \$4073 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1417 \$4075 \$1574 \$4074 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1418 \$4076 \$1574 \$4075 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1419 \$4077 \$1574 \$4076 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1420 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1421 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1422 \$4078 \$1574 \$3922 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1423 \$4079 \$1574 \$4078 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1424 \$4080 \$1574 \$4079 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1425 \$4081 \$1574 \$4080 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1426 \$4082 \$1574 \$4081 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1427 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1428 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1429 \$4083 \$1574 \$3927 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1430 \$4084 \$1574 \$4083 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1431 \$4085 \$1574 \$4084 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1432 \$4086 \$1574 \$4085 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1433 \$4087 \$1574 \$4086 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1434 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1435 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1436 \$4222 \$1573 \$3562 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1437 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1438 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1439 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1440 \$4224 \$1573 \$4223 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1441 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1442 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1443 \$4225 \$1573 \$3567 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1444 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1445 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1446 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1447 \$4227 \$1573 \$4226 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1448 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1449 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1450 \$4228 \$1573 \$3572 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1451 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1452 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1453 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1454 \$4230 \$1573 \$4229 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1455 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1456 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1457 \$4231 \$1574 \$3577 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1458 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1459 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1460 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1461 \$4232 \$1574 \$3582 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1462 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1463 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1464 \$4233 \$1574 \$3583 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1465 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1466 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1467 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1468 \$4234 \$1574 \$3588 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1469 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1470 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1471 \$4235 \$1574 \$3589 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1472 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1473 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1474 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1475 \$4236 \$1574 \$3594 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1476 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1477 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1478 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1479 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1480 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1481 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1482 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1483 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1484 \$4222 \$1573 \$4384 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1485 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1486 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1487 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1488 \$4224 \$1573 \$4385 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1489 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1490 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1491 \$4225 \$1573 \$4386 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1492 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1493 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1494 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1495 \$4227 \$1573 \$4387 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1496 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1497 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1498 \$4228 \$1573 \$4388 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1499 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1500 \$1573 \$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1501 AVDD|AVSS|VDD|VSS \$1573 \$1573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1502 \$4230 \$1573 \$4389 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1503 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1504 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1505 \$4231 \$1574 \$4390 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1506 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1507 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1508 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1509 \$4232 \$1574 \$32 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P
+ PS=5.3U PD=5.3U
M$1510 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1511 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1512 \$4233 \$1574 \$4391 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1513 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1514 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1515 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1516 \$4234 \$1574 \$33 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P
+ PS=5.3U PD=5.3U
M$1517 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1518 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1519 \$4235 \$1574 \$4392 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1520 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1521 AVDD|AVSS|VDD|VSS \$1574 \$1574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1522 \$1574 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1523 \$4236 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1524 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1525 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1526 \$4455 \$4383 \$1774 AVDD|AVSS|VDD|VSS pfet_03v3 L=6U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1527 AVDD|AVSS|VDD|VSS \$4383 \$4455 AVDD|AVSS|VDD|VSS pfet_03v3 L=6U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1528 \$4456 \$4383 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=6U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1529 \$1731 \$4383 \$4456 AVDD|AVSS|VDD|VSS pfet_03v3 L=6U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1530 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1531 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1532 \$4559 \$1573 \$4558 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1533 \$4560 \$1573 \$4559 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1534 \$4561 \$1573 \$4560 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1535 \$4562 \$1573 \$4561 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1536 \$4062 \$1573 \$4562 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1537 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1538 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1539 \$4564 \$1573 \$4563 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1540 \$4565 \$1573 \$4564 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1541 \$4566 \$1573 \$4565 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1542 \$4567 \$1573 \$4566 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1543 \$4067 \$1573 \$4567 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1544 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1545 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1546 \$4569 \$1573 \$4568 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1547 \$4570 \$1573 \$4569 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1548 \$4571 \$1573 \$4570 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1549 \$4572 \$1573 \$4571 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1550 \$4072 \$1573 \$4572 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1551 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1552 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1553 \$4574 \$1574 \$4573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1554 \$4575 \$1574 \$4574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1555 \$4576 \$1574 \$4575 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1556 \$4577 \$1574 \$4576 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1557 \$4077 \$1574 \$4577 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1558 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1559 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1560 \$4579 \$1574 \$4578 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1561 \$4580 \$1574 \$4579 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1562 \$4581 \$1574 \$4580 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1563 \$4582 \$1574 \$4581 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1564 \$4082 \$1574 \$4582 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1565 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1566 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1567 \$4584 \$1574 \$4583 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1568 \$4585 \$1574 \$4584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1569 \$4586 \$1574 \$4585 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1570 \$4587 \$1574 \$4586 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1571 \$4087 \$1574 \$4587 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1572 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1574 \$4638 \$4383 \$4383 AVDD|AVSS|VDD|VSS pfet_03v3 L=6U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1575 AVDD|AVSS|VDD|VSS \$4383 \$4638 AVDD|AVSS|VDD|VSS pfet_03v3 L=6U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1576 \$4639 \$4383 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=6U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1577 \$4383 \$4383 \$4639 AVDD|AVSS|VDD|VSS pfet_03v3 L=6U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1578 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1579 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1580 \$4741 \$1573 \$4558 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1581 \$4742 \$1573 \$4741 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1582 \$4743 \$1573 \$4742 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1583 \$4744 \$1573 \$4743 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1584 \$4745 \$1573 \$4744 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1585 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1586 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1587 \$4746 \$1573 \$4563 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1588 \$4747 \$1573 \$4746 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1589 \$4748 \$1573 \$4747 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1590 \$4749 \$1573 \$4748 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1591 \$4750 \$1573 \$4749 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1592 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1593 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1594 \$4751 \$1573 \$4568 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1595 \$4752 \$1573 \$4751 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1596 \$4753 \$1573 \$4752 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1597 \$4754 \$1573 \$4753 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1598 \$4755 \$1573 \$4754 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1599 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1600 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1601 \$4756 \$1574 \$4573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1602 \$4757 \$1574 \$4756 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1603 \$4758 \$1574 \$4757 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1604 \$4759 \$1574 \$4758 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1605 \$4760 \$1574 \$4759 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1606 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1607 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1608 \$4761 \$1574 \$4578 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1609 \$4762 \$1574 \$4761 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1610 \$4763 \$1574 \$4762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1611 \$4764 \$1574 \$4763 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1612 \$4765 \$1574 \$4764 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1613 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1614 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1615 \$4766 \$1574 \$4583 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1616 \$4767 \$1574 \$4766 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1617 \$4768 \$1574 \$4767 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1618 \$4769 \$1574 \$4768 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1619 \$4770 \$1574 \$4769 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1620 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1621 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1622 \$4812 \$4383 \$1731 AVDD|AVSS|VDD|VSS pfet_03v3 L=6U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1623 AVDD|AVSS|VDD|VSS \$4383 \$4812 AVDD|AVSS|VDD|VSS pfet_03v3 L=6U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1624 \$4813 \$4383 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=6U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1625 \$1774 \$4383 \$4813 AVDD|AVSS|VDD|VSS pfet_03v3 L=6U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1626 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1627 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1628 \$4912 \$1573 \$6255 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1629 \$4913 \$1573 \$4912 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1630 \$4914 \$1573 \$4913 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1631 \$4915 \$1573 \$4914 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1632 \$4745 \$1573 \$4915 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1633 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1634 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1635 \$4916 \$1573 \$6256 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1636 \$4917 \$1573 \$4916 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1637 \$4918 \$1573 \$4917 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1638 \$4919 \$1573 \$4918 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1639 \$4750 \$1573 \$4919 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1640 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1641 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1642 \$4920 \$1573 \$6257 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1643 \$4921 \$1573 \$4920 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1644 \$4922 \$1573 \$4921 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1645 \$4923 \$1573 \$4922 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1646 \$4755 \$1573 \$4923 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1647 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1648 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1649 \$4924 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1650 \$4925 \$1574 \$4924 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1651 \$4926 \$1574 \$4925 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1652 \$4927 \$1574 \$4926 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1653 \$4760 \$1574 \$4927 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1654 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1655 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1656 \$4928 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1657 \$4929 \$1574 \$4928 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1658 \$4930 \$1574 \$4929 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1659 \$4931 \$1574 \$4930 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1660 \$4765 \$1574 \$4931 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1661 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1662 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1663 \$4932 \$1574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1664 \$4933 \$1574 \$4932 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1665 \$4934 \$1574 \$4933 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1666 \$4935 \$1574 \$4934 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1667 \$4770 \$1574 \$4935 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1668 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1669 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1670 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1671 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1672 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1673 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1674 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1675 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1676 \$5053 \$1573 \$4384 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1677 \$5054 \$1573 \$5053 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1678 \$5055 \$1573 \$5054 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1679 \$5056 \$1573 \$5055 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1680 \$4385 \$1573 \$5056 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1681 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1682 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1683 \$5057 \$1573 \$4386 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1684 \$5058 \$1573 \$5057 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1685 \$5059 \$1573 \$5058 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1686 \$5060 \$1573 \$5059 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1687 \$4387 \$1573 \$5060 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1688 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1689 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1690 \$5061 \$1573 \$4388 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1691 \$5062 \$1573 \$5061 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1692 \$5063 \$1573 \$5062 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1693 \$5064 \$1573 \$5063 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1694 \$4389 \$1573 \$5064 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1695 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1696 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1697 \$5065 \$1574 \$4390 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1698 \$5066 \$1574 \$5065 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1699 \$5067 \$1574 \$5066 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1700 \$5068 \$1574 \$5067 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1701 AVDD|AVSS|VDD|VSS \$1574 \$5068 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1702 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1703 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1704 \$5069 \$1574 \$4391 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1705 \$5070 \$1574 \$5069 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1706 \$5071 \$1574 \$5070 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1707 \$5072 \$1574 \$5071 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1708 AVDD|AVSS|VDD|VSS \$1574 \$5072 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1709 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1710 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1711 \$5073 \$1574 \$4392 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=1.3P PS=5.3U PD=5.3U
M$1712 \$5074 \$1574 \$5073 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1713 \$5075 \$1574 \$5074 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$1714 \$5076 \$1574 \$5075 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1715 AVDD|AVSS|VDD|VSS \$1574 \$5076 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1716 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1717 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1718 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1719 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1720 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1721 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1722 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1723 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1724 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1725 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1726 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1727 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1728 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1729 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1730 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1731 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1732 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1733 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1734 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1735 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1736 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1737 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1738 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1739 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1740 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1741 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1742 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1743 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1744 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1745 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1746 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1747 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1748 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1749 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1750 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1751 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1752 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1753 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1754 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1755 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1756 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1757 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1758 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1759 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1760 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1761 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1762 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1763 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1764 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1765 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1766 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1767 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1768 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1769 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1770 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1771 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1772 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1773 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1774 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1775 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1776 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1777 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1778 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1779 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1780 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1781 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1782 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1783 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1784 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1785 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1786 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1787 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1788 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1789 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1790 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1791 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1792 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1793 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1794 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1795 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1796 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1797 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1798 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1799 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1800 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1801 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1802 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1803 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1804 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1805 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1806 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1807 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1808 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1809 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1810 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1811 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1812 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1813 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1814 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1815 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1816 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1817 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1818 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1819 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1820 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1821 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1822 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1823 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1824 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1825 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1826 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1827 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1828 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1829 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1830 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1831 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1832 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1833 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1834 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1835 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1836 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1837 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1838 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1839 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1840 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1841 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1842 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1843 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1844 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1845 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1846 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1847 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1848 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1849 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1850 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1851 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1852 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1853 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1854 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1855 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1856 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1857 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1858 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1859 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1860 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1861 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1862 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1863 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1864 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1865 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1866 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1867 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1868 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1869 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1870 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1871 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1872 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1873 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1874 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1875 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1876 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1877 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1878 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1879 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1880 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1881 \$6116 \$5372 \$5372 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1882 AVDD|AVSS|VDD|VSS \$5372 \$6116 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1883 \$6117 \$5372 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1884 \$5271 \$5372 \$6117 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1885 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1886 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1887 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1888 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1889 \$6118 \$6150 A1|VN AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1890 \$5375 \$6150 \$6118 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1891 \$6119 \$6150 \$5482 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1892 \$6120 \$6150 \$6119 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1893 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1894 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1895 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1896 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1897 \$6121 \$5472 \$5473 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1898 \$4223 \$5472 \$6121 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1899 \$6122 \$6255 \$4223 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1900 \$6150 \$6255 \$6122 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1901 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1902 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1903 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1904 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1905 \$6123 \$5380 \$5380 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1906 AVDD|AVSS|VDD|VSS \$5380 \$6123 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1907 \$6124 \$5380 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1908 \$5272 \$5380 \$6124 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1909 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1910 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1911 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1912 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1913 \$6125 \$6151 \$6120 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1914 \$5383 \$6151 \$6125 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1915 \$6126 \$6151 \$5483 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1916 \$6127 \$6151 \$6126 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1917 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1918 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1919 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1920 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1921 \$6128 \$5474 \$5475 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1922 \$4226 \$5474 \$6128 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1923 \$6129 \$6256 \$4226 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1924 \$6151 \$6256 \$6129 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1925 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1926 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1927 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1928 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1929 \$6130 \$5388 \$5388 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1930 AVDD|AVSS|VDD|VSS \$5388 \$6130 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1931 \$6131 \$5388 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1932 \$5273 \$5388 \$6131 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1933 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1934 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1935 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1936 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1937 \$6132 \$6152 \$6127 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1938 \$5391 \$6152 \$6132 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1939 \$6133 \$6152 \$5484 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1940 \$6134 \$6152 \$6133 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1941 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1942 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1943 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1944 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1945 \$6135 \$5476 \$5477 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1946 \$4229 \$5476 \$6135 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1947 \$6136 \$6257 \$4229 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1948 \$6152 \$6257 \$6136 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1949 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1950 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1951 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1952 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1953 \$6137 \$5396 \$5396 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1954 AVDD|AVSS|VDD|VSS \$5396 \$6137 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1955 \$6138 \$5396 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1956 \$5274 \$5396 \$6138 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1957 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1958 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1959 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1960 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1961 \$6139 \$6153 \$6134 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1962 \$5399 \$6153 \$6139 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1963 \$6140 \$6153 \$5485 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1964 \$6141 \$6153 \$6140 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1965 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1966 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1967 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1968 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1969 \$6142 \$5478 \$5479 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1970 \$2148 \$5478 \$6142 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1971 \$6143 \$6258 \$2148 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1972 \$6153 \$6258 \$6143 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1973 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1974 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1975 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1976 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1977 \$6144 \$5404 \$5404 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1978 AVDD|AVSS|VDD|VSS \$5404 \$6144 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1979 \$6145 \$5404 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1980 \$5275 \$5404 \$6145 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1981 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1982 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1983 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1984 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1985 \$6146 \$6154 \$6141 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1986 \$5407 \$6154 \$6146 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1987 \$6147 \$6154 \$5486 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1988 B1|VOUT \$6154 \$6147 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1989 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1990 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1991 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1992 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1993 \$6148 \$5480 \$5481 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1994 \$2151 \$5480 \$6148 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1995 \$6149 \$6259 \$2151 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$1996 \$6154 \$6259 \$6149 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$1997 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1998 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1999 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2000 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2001 \$6275 \$5372 \$5271 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2002 AVDD|AVSS|VDD|VSS \$5372 \$6275 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2003 \$6276 \$5372 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2004 \$5372 \$5372 \$6276 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2005 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2006 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2007 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2008 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2009 \$6277 \$6150 \$6255 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2010 AVDD|AVSS|VDD|VSS \$6150 \$6277 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2011 \$6278 \$6150 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2012 \$6255 \$6150 \$6278 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2013 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2014 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2015 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2016 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2017 \$6279 \$6255 \$6150 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2018 \$4223 \$6255 \$6279 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2019 \$6280 \$5472 \$4223 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2020 \$5473 \$5472 \$6280 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2021 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2022 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2023 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2024 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2025 \$6281 \$5380 \$5272 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2026 AVDD|AVSS|VDD|VSS \$5380 \$6281 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2027 \$6282 \$5380 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2028 \$5380 \$5380 \$6282 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2029 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2030 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2031 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2032 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2033 \$6283 \$6151 \$6256 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2034 AVDD|AVSS|VDD|VSS \$6151 \$6283 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2035 \$6284 \$6151 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2036 \$6256 \$6151 \$6284 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2037 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2038 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2039 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2040 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2041 \$6285 \$6256 \$6151 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2042 \$4226 \$6256 \$6285 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2043 \$6286 \$5474 \$4226 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2044 \$5475 \$5474 \$6286 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2045 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2046 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2047 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2048 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2049 \$6287 \$5388 \$5273 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2050 AVDD|AVSS|VDD|VSS \$5388 \$6287 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2051 \$6288 \$5388 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2052 \$5388 \$5388 \$6288 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2053 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2054 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2055 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2056 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2057 \$6289 \$6152 \$6257 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2058 AVDD|AVSS|VDD|VSS \$6152 \$6289 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2059 \$6290 \$6152 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2060 \$6257 \$6152 \$6290 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2061 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2062 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2063 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2064 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2065 \$6291 \$6257 \$6152 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2066 \$4229 \$6257 \$6291 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2067 \$6292 \$5476 \$4229 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2068 \$5477 \$5476 \$6292 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2069 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2070 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2071 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2072 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2073 \$6293 \$5396 \$5274 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2074 AVDD|AVSS|VDD|VSS \$5396 \$6293 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2075 \$6294 \$5396 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2076 \$5396 \$5396 \$6294 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2077 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2078 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2079 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2080 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2081 \$6295 \$6153 \$6258 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2082 AVDD|AVSS|VDD|VSS \$6153 \$6295 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2083 \$6296 \$6153 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2084 \$6258 \$6153 \$6296 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2085 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2086 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2087 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2088 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2089 \$6297 \$6258 \$6153 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2090 \$2148 \$6258 \$6297 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2091 \$6298 \$5478 \$2148 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2092 \$5479 \$5478 \$6298 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2093 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2094 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2095 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2096 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2097 \$6299 \$5404 \$5275 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2098 AVDD|AVSS|VDD|VSS \$5404 \$6299 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2099 \$6300 \$5404 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2100 \$5404 \$5404 \$6300 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2101 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2102 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2103 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2104 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2105 \$6301 \$6154 \$6259 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2106 AVDD|AVSS|VDD|VSS \$6154 \$6301 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2107 \$6302 \$6154 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2108 \$6259 \$6154 \$6302 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2109 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2110 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2111 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2112 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2113 \$6303 \$6259 \$6154 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2114 \$2151 \$6259 \$6303 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2115 \$6304 \$5480 \$2151 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2116 \$5481 \$5480 \$6304 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2117 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2118 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2119 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2120 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2121 \$6411 \$5372 \$5372 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2122 AVDD|AVSS|VDD|VSS \$5372 \$6411 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2123 \$6412 \$5372 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2124 \$5271 \$5372 \$6412 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2125 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2126 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2127 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2128 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2129 \$6413 \$6150 \$6255 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2130 AVDD|AVSS|VDD|VSS \$6150 \$6413 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2131 \$6414 \$6150 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2132 \$6255 \$6150 \$6414 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2133 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2134 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2135 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2136 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2137 \$6415 \$5472 \$5473 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2138 \$4223 \$5472 \$6415 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2139 \$6416 \$6255 \$4223 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2140 \$6150 \$6255 \$6416 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2141 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2142 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2143 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2144 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2145 \$6417 \$5380 \$5380 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2146 AVDD|AVSS|VDD|VSS \$5380 \$6417 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2147 \$6418 \$5380 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2148 \$5272 \$5380 \$6418 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2149 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2150 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2151 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2152 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2153 \$6419 \$6151 \$6256 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2154 AVDD|AVSS|VDD|VSS \$6151 \$6419 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2155 \$6420 \$6151 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2156 \$6256 \$6151 \$6420 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2157 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2158 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2159 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2160 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2161 \$6421 \$5474 \$5475 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2162 \$4226 \$5474 \$6421 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2163 \$6422 \$6256 \$4226 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2164 \$6151 \$6256 \$6422 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2165 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2166 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2167 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2168 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2169 \$6423 \$5388 \$5388 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2170 AVDD|AVSS|VDD|VSS \$5388 \$6423 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2171 \$6424 \$5388 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2172 \$5273 \$5388 \$6424 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2173 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2174 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2175 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2176 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2177 \$6425 \$6152 \$6257 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2178 AVDD|AVSS|VDD|VSS \$6152 \$6425 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2179 \$6426 \$6152 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2180 \$6257 \$6152 \$6426 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2181 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2182 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2183 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2184 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2185 \$6427 \$5476 \$5477 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2186 \$4229 \$5476 \$6427 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2187 \$6428 \$6257 \$4229 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2188 \$6152 \$6257 \$6428 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2189 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2190 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2191 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2192 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2193 \$6429 \$5396 \$5396 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2194 AVDD|AVSS|VDD|VSS \$5396 \$6429 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2195 \$6430 \$5396 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2196 \$5274 \$5396 \$6430 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2197 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2198 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2199 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2200 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2201 \$6431 \$6153 \$6258 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2202 AVDD|AVSS|VDD|VSS \$6153 \$6431 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2203 \$6432 \$6153 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2204 \$6258 \$6153 \$6432 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2205 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2206 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2207 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2208 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2209 \$6433 \$5478 \$5479 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2210 \$2148 \$5478 \$6433 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2211 \$6434 \$6258 \$2148 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2212 \$6153 \$6258 \$6434 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2213 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2214 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2215 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2216 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2217 \$6435 \$5404 \$5404 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2218 AVDD|AVSS|VDD|VSS \$5404 \$6435 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2219 \$6436 \$5404 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2220 \$5275 \$5404 \$6436 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2221 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2222 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2223 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2224 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2225 \$6437 \$6154 \$6259 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2226 AVDD|AVSS|VDD|VSS \$6154 \$6437 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2227 \$6438 \$6154 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2228 \$6259 \$6154 \$6438 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2229 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2230 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2231 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2232 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2233 \$6439 \$5480 \$5481 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2234 \$2151 \$5480 \$6439 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2235 \$6440 \$6259 \$2151 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2236 \$6154 \$6259 \$6440 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2237 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2238 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2239 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2240 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2241 \$6571 \$5372 \$5271 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2242 AVDD|AVSS|VDD|VSS \$5372 \$6571 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2243 \$6572 \$5372 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2244 \$5372 \$5372 \$6572 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2245 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2246 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2247 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2248 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2249 \$6573 \$6150 \$6120 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2250 \$5482 \$6150 \$6573 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2251 \$6574 \$6150 \$5375 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2252 A1|VN \$6150 \$6574 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2253 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2254 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2255 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2256 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2257 \$6575 \$6255 \$6150 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2258 \$4223 \$6255 \$6575 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2259 \$6576 \$5472 \$4223 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2260 \$5473 \$5472 \$6576 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2261 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2263 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2264 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2265 \$6577 \$5380 \$5272 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2266 AVDD|AVSS|VDD|VSS \$5380 \$6577 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2267 \$6578 \$5380 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2268 \$5380 \$5380 \$6578 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2269 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2270 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2271 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2272 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2273 \$6579 \$6151 \$6127 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2274 \$5483 \$6151 \$6579 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2275 \$6580 \$6151 \$5383 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2276 \$6120 \$6151 \$6580 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2277 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2278 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2279 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2280 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2281 \$6581 \$6256 \$6151 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2282 \$4226 \$6256 \$6581 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2283 \$6582 \$5474 \$4226 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2284 \$5475 \$5474 \$6582 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2285 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2286 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2287 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2288 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2289 \$6583 \$5388 \$5273 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2290 AVDD|AVSS|VDD|VSS \$5388 \$6583 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2291 \$6584 \$5388 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2292 \$5388 \$5388 \$6584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2293 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2294 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2295 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2296 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2297 \$6585 \$6152 \$6134 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2298 \$5484 \$6152 \$6585 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2299 \$6586 \$6152 \$5391 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2300 \$6127 \$6152 \$6586 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2301 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2302 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2303 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2304 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2305 \$6587 \$6257 \$6152 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2306 \$4229 \$6257 \$6587 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2307 \$6588 \$5476 \$4229 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2308 \$5477 \$5476 \$6588 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2309 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2310 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2311 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2312 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2313 \$6589 \$5396 \$5274 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2314 AVDD|AVSS|VDD|VSS \$5396 \$6589 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2315 \$6590 \$5396 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2316 \$5396 \$5396 \$6590 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2317 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2318 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2319 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2320 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2321 \$6591 \$6153 \$6141 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2322 \$5485 \$6153 \$6591 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2323 \$6592 \$6153 \$5399 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2324 \$6134 \$6153 \$6592 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2325 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2326 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2327 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2328 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2329 \$6593 \$6258 \$6153 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2330 \$2148 \$6258 \$6593 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2331 \$6594 \$5478 \$2148 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2332 \$5479 \$5478 \$6594 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2333 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2334 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2335 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2336 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2337 \$6595 \$5404 \$5275 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2338 AVDD|AVSS|VDD|VSS \$5404 \$6595 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2339 \$6596 \$5404 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2340 \$5404 \$5404 \$6596 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2341 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2342 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2343 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2344 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2345 \$6597 \$6154 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2346 \$5486 \$6154 \$6597 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2347 \$6598 \$6154 \$5407 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2348 \$6141 \$6154 \$6598 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2349 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2350 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2351 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2352 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2353 \$6599 \$6259 \$6154 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2354 \$2151 \$6259 \$6599 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2355 \$6600 \$5480 \$2151 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2356 \$5481 \$5480 \$6600 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2357 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2358 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2359 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2360 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2361 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2362 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2363 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2364 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2365 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2366 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2367 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2368 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2369 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2370 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2371 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2372 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2373 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2374 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2375 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2376 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2377 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2378 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2379 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2380 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2381 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2382 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2383 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2384 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2385 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2386 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2387 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2388 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2389 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2390 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2391 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2392 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2393 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2394 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2395 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2396 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2397 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2398 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2399 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2400 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2401 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2402 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2403 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2404 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2405 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2406 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2407 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2408 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2409 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2410 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2411 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2412 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2413 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2414 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2415 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2416 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2417 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2418 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2419 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2420 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2421 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2422 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2423 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2424 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2425 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2426 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2427 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2428 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2429 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2430 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2431 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2432 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2433 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2434 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2435 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2436 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2437 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2438 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2439 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2440 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2441 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2442 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2443 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2444 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2445 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2446 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2447 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2448 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2449 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2450 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2451 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2452 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2453 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2454 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2455 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2456 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2457 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2458 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2459 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2460 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2461 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2462 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2463 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2464 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2465 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2466 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2467 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2468 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2469 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2470 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2471 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2472 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2473 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2474 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2475 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2476 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2477 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2478 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2479 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2480 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2481 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2482 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2483 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2484 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2485 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2486 AVDD|AVSS|VDD|VSS IREF \$6812 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2487 \$6812 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2488 AVDD|AVSS|VDD|VSS IREF \$6812 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2489 \$6812 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2490 AVDD|AVSS|VDD|VSS IREF \$6843 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2491 \$6843 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2492 AVDD|AVSS|VDD|VSS IREF \$6843 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2493 \$6843 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2494 AVDD|AVSS|VDD|VSS IREF IREF AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2495 IREF IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2496 AVDD|AVSS|VDD|VSS IREF IREF AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2497 IREF IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2498 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2499 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2500 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2501 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2502 AVDD|AVSS|VDD|VSS IREF IREF AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2503 IREF IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2504 AVDD|AVSS|VDD|VSS IREF IREF AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2505 IREF IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2506 AVDD|AVSS|VDD|VSS IREF \$6843 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2507 \$6843 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2508 AVDD|AVSS|VDD|VSS IREF \$6843 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2509 \$6843 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2510 AVDD|AVSS|VDD|VSS IREF \$6812 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2511 \$6812 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2512 AVDD|AVSS|VDD|VSS IREF \$6812 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2513 \$6812 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2514 AVDD|AVSS|VDD|VSS IREF IREF AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2515 IREF IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2516 AVDD|AVSS|VDD|VSS IREF IREF AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2517 AVDD|AVSS|VDD|VSS IREF \$6843 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2518 \$6843 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2519 AVDD|AVSS|VDD|VSS IREF \$6843 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2520 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2521 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2522 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2523 \$6843 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2524 AVDD|AVSS|VDD|VSS IREF \$6843 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2525 \$6843 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2526 \$6812 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2527 AVDD|AVSS|VDD|VSS IREF \$6812 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2528 \$6812 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2529 AVDD|AVSS|VDD|VSS IREF \$6812 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2530 \$6812 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2531 AVDD|AVSS|VDD|VSS IREF \$6812 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2532 AVDD|AVSS|VDD|VSS IREF IREF AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2533 IREF IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2534 AVDD|AVSS|VDD|VSS IREF IREF AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2535 AVDD|AVSS|VDD|VSS IREF IREF AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2536 IREF IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2537 AVDD|AVSS|VDD|VSS IREF IREF AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2538 IREF IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2539 AVDD|AVSS|VDD|VSS IREF \$6843 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2540 \$6843 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2541 AVDD|AVSS|VDD|VSS IREF \$6843 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2542 \$6843 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2543 AVDD|AVSS|VDD|VSS IREF \$6843 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2544 \$6843 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2545 AVDD|AVSS|VDD|VSS IREF \$6843 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2546 \$6843 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2547 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2548 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2549 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2550 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2551 AVDD|AVSS|VDD|VSS IREF \$6812 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2552 \$6812 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2553 AVDD|AVSS|VDD|VSS IREF \$6812 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2554 \$6812 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2555 AVDD|AVSS|VDD|VSS IREF IREF AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2556 IREF IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2557 AVDD|AVSS|VDD|VSS IREF IREF AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2558 IREF IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2559 AVDD|AVSS|VDD|VSS IREF \$6812 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2560 \$6812 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2561 AVDD|AVSS|VDD|VSS IREF \$6812 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2562 \$6812 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2563 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2564 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2565 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2566 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2567 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2568 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2569 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2570 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2571 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2572 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2575 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2576 \$10774 \$6797 \$10096 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=1.2U AS=0.78P
+ AD=0.504P PS=3.7U PD=2.04U
M$2577 \$10775 \$6797 \$10774 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=1.2U AS=0.504P
+ AD=0.504P PS=2.04U PD=2.04U
M$2578 \$10776 \$6797 \$10775 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=1.2U AS=0.504P
+ AD=0.78P PS=2.04U PD=3.7U
M$2579 \$11315 \$6797 \$11314 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=1.2U AS=0.78P
+ AD=0.504P PS=3.7U PD=2.04U
M$2580 \$11316 \$6797 \$11315 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=1.2U AS=0.504P
+ AD=0.504P PS=2.04U PD=2.04U
M$2581 \$10776 \$6797 \$11316 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=1.2U AS=0.504P
+ AD=0.78P PS=2.04U PD=3.7U
M$2582 \$10097 \$6797 \$10096 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=1.2U AS=0.78P
+ AD=0.504P PS=3.7U PD=2.04U
M$2583 \$10098 \$6797 \$10097 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=1.2U AS=0.504P
+ AD=0.504P PS=2.04U PD=2.04U
M$2584 AVDD|AVSS|VDD|VSS \$6797 \$10098 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=1.2U
+ AS=0.504P AD=0.78P PS=2.04U PD=3.7U
M$2585 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P PS=3.7U PD=2.04U
M$2586 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P PS=2.04U PD=2.04U
M$2587 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P PS=2.04U PD=3.7U
M$2588 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P PS=3.7U PD=2.04U
M$2589 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P PS=2.04U PD=2.04U
M$2590 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P PS=2.04U PD=3.7U
M$2591 \$11850 \$6797 \$11314 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=1.2U AS=0.78P
+ AD=0.504P PS=3.7U PD=2.04U
M$2592 \$11851 \$6797 \$11850 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=1.2U AS=0.504P
+ AD=0.504P PS=2.04U PD=2.04U
M$2593 \$11852 \$6797 \$11851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=1.2U AS=0.504P
+ AD=0.78P PS=2.04U PD=3.7U
M$2594 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2595 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2596 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2597 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2598 \$6797 \$6797 \$11852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=1.2U AS=0.78P
+ AD=0.78P PS=3.7U PD=3.7U
M$2599 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2600 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2601 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2602 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2603 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2604 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2605 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2606 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2607 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2608 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2609 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2610 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2611 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2612 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2613 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2614 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2615 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2616 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2617 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2618 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2619 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2620 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2621 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2622 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2623 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2624 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2625 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2626 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2627 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2628 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2629 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2630 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2631 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2632 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2633 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2634 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2635 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2636 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2637 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2638 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2639 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2640 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2641 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2642 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2643 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2644 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2645 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2646 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2647 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2648 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2649 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2650 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2651 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2652 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2653 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2654 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2655 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2656 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2657 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2658 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2659 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2660 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2661 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2662 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2663 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2664 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2665 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2666 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2667 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2668 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2669 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2670 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2671 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2672 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2673 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2674 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2675 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2676 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2677 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2678 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2679 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2680 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2681 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2682 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2683 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2684 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2685 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2686 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2687 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2688 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2689 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2690 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2691 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2692 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2693 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2694 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2695 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2696 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2697 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2698 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2699 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2700 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2701 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2702 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2703 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2704 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2705 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2706 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2707 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2708 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2709 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2710 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2711 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2712 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2713 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2714 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2715 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2716 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2717 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2718 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2719 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2720 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2721 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2722 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2723 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2724 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2725 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2726 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2727 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2728 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2729 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2730 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2731 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2732 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2733 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2734 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2735 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2736 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2737 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2738 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2739 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2740 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2741 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2742 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2743 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2744 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2745 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2746 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2747 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2748 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2749 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2750 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2751 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2752 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2753 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2754 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2755 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2756 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2757 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2758 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2759 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2760 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2761 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2762 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2763 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2764 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2765 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2766 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2767 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2768 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2769 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2770 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2771 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2772 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2773 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2774 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2775 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2776 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2777 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2778 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2779 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2780 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2781 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2782 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2783 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2784 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2785 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2786 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2787 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2788 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2789 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2790 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2791 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2792 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2793 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2794 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2795 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2796 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2797 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2798 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2799 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2800 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2801 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2802 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2803 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2804 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2805 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2806 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2807 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2808 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2809 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2810 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2811 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2812 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2813 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2814 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2815 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2816 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2817 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2818 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2819 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2820 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2821 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2822 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2823 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2824 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2825 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2826 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2827 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2828 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2829 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2830 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2831 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2832 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2833 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2834 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2835 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2836 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2837 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2838 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2839 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2840 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2841 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2842 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2843 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2844 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2845 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2846 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2847 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2848 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2849 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2850 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2851 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2852 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2853 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2854 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2855 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2856 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2857 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2858 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2859 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2860 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2861 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2862 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2863 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2864 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2865 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2866 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2867 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2868 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2869 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2870 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2871 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2872 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2873 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2874 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2875 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2876 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2877 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2878 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2879 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2880 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2881 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2882 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2883 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2884 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2885 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2886 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2887 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2888 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2889 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2890 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2891 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2892 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2893 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2894 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2895 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2896 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2897 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2898 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2899 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2900 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2901 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2902 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2903 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2904 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2905 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2906 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2907 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2908 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2909 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2910 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2911 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2912 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2913 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2914 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2915 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2916 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2917 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2918 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2919 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2920 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2921 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2922 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2923 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2924 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2925 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2926 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2927 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2928 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2929 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2930 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2931 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2932 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2933 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2934 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2935 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2936 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2937 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2938 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2939 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2940 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2941 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2942 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2943 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2944 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2945 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2946 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2947 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2948 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2949 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2950 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2951 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2952 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2953 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2954 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2955 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2956 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2957 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2958 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2959 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2960 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2961 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2962 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2963 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2964 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2965 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2966 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2967 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2968 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2969 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2970 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2971 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2972 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2973 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2974 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2975 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2976 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2977 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2978 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2979 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2980 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2981 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2982 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2983 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2984 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2985 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2986 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2987 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2988 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$2989 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2990 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$2991 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2992 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2993 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2994 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2995 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2996 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2997 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$2998 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$2999 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3000 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3001 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3002 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3003 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3004 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$3005 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3006 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3007 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3008 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3009 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3010 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3011 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3012 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3013 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3014 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3015 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3016 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3017 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3018 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3019 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3020 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3021 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3022 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3023 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3024 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3025 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3026 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3027 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3028 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3029 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3030 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3031 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3032 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3033 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3034 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3035 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3036 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3037 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3038 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3039 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3040 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$3041 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3042 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3043 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3044 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3045 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3046 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3047 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3048 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3049 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3050 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3051 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3052 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3053 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$3054 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3055 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3056 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3057 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3058 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3059 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3060 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3061 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3062 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3063 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3064 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3065 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3066 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3067 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3068 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3069 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3070 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3071 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3072 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3073 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3074 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3075 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3076 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3077 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3078 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3079 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3080 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3081 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3082 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3083 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3084 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3085 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3086 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3087 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3088 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3089 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3090 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3091 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3092 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$3093 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3094 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3095 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3096 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3097 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3098 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3099 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3100 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3101 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3102 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3103 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3104 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3105 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$3106 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3107 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3108 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3109 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3110 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3111 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3112 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3113 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3114 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3115 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3116 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3117 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3118 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3119 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3120 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3121 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3122 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3123 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3124 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3125 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3126 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3127 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3128 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3129 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3130 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3131 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3132 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3133 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3134 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3135 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3136 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3137 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3138 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3139 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3140 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$3141 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3142 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3143 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3144 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3145 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3146 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3147 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$3148 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3149 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3150 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3151 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3152 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3153 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$3154 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3155 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3156 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3157 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3158 \$19851 A1|VN \$6762 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3159 \$6762 A1|VN \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3160 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P
+ PS=5.3U PD=2.84U
M$3161 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3162 \$19851 VP \$6793 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3163 \$6793 VP \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3164 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3165 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3166 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3167 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3168 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3169 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3170 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3171 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3172 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3173 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3174 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3175 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3176 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3177 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3178 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3179 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3180 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3181 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3182 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3183 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3184 \$19584 \$6797 B1|VOUT AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3185 B1|VOUT \$6797 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3186 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=1.3P
+ AD=0.84P PS=5.3U PD=2.84U
M$3187 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3188 \$19852 \$6797 \$12262 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=0.84P PS=2.84U PD=2.84U
M$3189 \$12262 \$6797 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U AS=0.84P
+ AD=1.3P PS=2.84U PD=5.3U
M$3190 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3191 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3192 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3193 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3194 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3195 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3196 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3197 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3198 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3199 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3200 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3201 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3202 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3203 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3204 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3205 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3206 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3207 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3208 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3209 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3210 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3211 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3212 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3213 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3214 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3215 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3216 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3217 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3218 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3219 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3220 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3221 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3222 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3223 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3224 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3225 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3226 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3227 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3228 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3229 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3230 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3231 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3232 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3233 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3234 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3235 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3236 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3237 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3238 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3239 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3240 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3241 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3242 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3243 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3244 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3245 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3246 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3247 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3248 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3249 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3250 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3251 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3252 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3253 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3254 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3255 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3256 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3257 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3258 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3259 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3260 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3261 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3263 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3264 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3265 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3266 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3267 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3268 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3269 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3270 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3271 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3272 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3273 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3274 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3275 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3276 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3277 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3278 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3279 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3280 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3281 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3282 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3283 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3284 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3285 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3286 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3287 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3288 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3289 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3290 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3291 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3292 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3293 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3294 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3295 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3296 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3297 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3298 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3299 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3300 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3301 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3302 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3303 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3304 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3305 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3306 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3307 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3308 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3309 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3310 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3311 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3312 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3313 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3314 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3315 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3316 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3317 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3318 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3319 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3320 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3321 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3322 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3323 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3324 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3325 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3326 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3327 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3328 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3329 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3330 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3331 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3332 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3333 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3334 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3335 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3336 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3337 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3338 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3339 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3340 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3341 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3342 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3343 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3344 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3345 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3346 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3347 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3348 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3349 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3350 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3351 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3352 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3353 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3354 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3355 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3356 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3357 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3358 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3359 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3360 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3361 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3362 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3363 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3364 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3365 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3366 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3367 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3368 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3369 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3370 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3371 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3372 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3373 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3374 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3375 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3376 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3377 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3378 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3379 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3380 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3381 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3382 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3383 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3384 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3385 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3386 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3387 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3388 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3389 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3390 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3391 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3392 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3393 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3394 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3395 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3396 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3397 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3398 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3399 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3400 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3401 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3402 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3403 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3404 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3405 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3406 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3407 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3408 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3409 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3410 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3411 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3412 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3413 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3414 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3415 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3416 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3417 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3418 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3419 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3420 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3421 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3422 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3423 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3424 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3425 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3426 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3427 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3428 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3429 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3430 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3431 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3432 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3433 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3434 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3435 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3436 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3437 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3438 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3439 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3440 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3441 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3442 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3443 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3444 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3445 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3446 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3447 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3448 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3449 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3450 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3451 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3452 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3453 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3454 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3455 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3456 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3457 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3458 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3459 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3460 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3461 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3462 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3463 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3464 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3465 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3466 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3467 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3468 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3469 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3470 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3471 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3472 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3473 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3474 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3475 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3476 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3477 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3478 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3479 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3480 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3481 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3482 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3483 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3484 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3485 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3486 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3487 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3488 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3489 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3490 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3491 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3492 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3493 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3494 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3495 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3496 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3497 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3498 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3499 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3500 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3501 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3502 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3503 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3504 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3505 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3506 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3507 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3508 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3509 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3510 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3511 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3512 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3513 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3514 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3515 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3516 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3517 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3518 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3519 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3520 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3521 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3522 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3523 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3524 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3525 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3526 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3527 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3528 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3529 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3530 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3531 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3532 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3533 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3534 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3535 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3536 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3537 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3538 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3539 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3540 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3541 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3542 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3543 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3544 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3545 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3546 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3547 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3548 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3549 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3550 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3551 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3552 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3553 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3554 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3555 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3556 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3557 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3558 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3559 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3560 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3561 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3562 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3563 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3564 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3565 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3566 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3567 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3568 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3569 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3570 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3571 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3572 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3575 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3576 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3577 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3578 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3579 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3580 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3581 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3582 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3583 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3584 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3585 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3586 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3587 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3588 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3589 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3590 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3591 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3592 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3593 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3594 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3595 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3596 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3597 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3598 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3599 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3600 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3601 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3602 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3603 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3604 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3605 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3606 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3607 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3608 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3609 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3610 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3611 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3612 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3613 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3614 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3615 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3616 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3617 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3618 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3619 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3620 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3621 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3622 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3623 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3624 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3625 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3626 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3627 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3628 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3629 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3630 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3631 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3632 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3633 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3634 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3635 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3636 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3637 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3638 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3639 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3640 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3641 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3642 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3643 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3644 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3645 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3646 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3647 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3648 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3649 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3650 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3651 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3652 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3653 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3654 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3655 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3656 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3657 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3658 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3659 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3660 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3661 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3662 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3663 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3664 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3665 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3666 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3667 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3668 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3669 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3670 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3671 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3672 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3673 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3674 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3675 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3676 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3677 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3678 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3679 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3680 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3681 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3682 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3683 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3684 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3685 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3686 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3687 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3688 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3689 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3690 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3691 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3692 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3693 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3694 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3695 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3696 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3697 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3698 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3699 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3700 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3701 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3702 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3703 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3704 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3705 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3706 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3707 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3708 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3709 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3710 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3711 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3712 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3713 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3714 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3715 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3716 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3717 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3718 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3719 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3720 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3721 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3722 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3723 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3724 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3725 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3726 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3727 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3728 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3729 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3730 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3731 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3732 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3733 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3734 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3735 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3736 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3737 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3738 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3739 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3740 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3741 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3742 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3743 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3744 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3745 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3746 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3747 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3748 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3749 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3750 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3751 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3752 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3753 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3754 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3755 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3756 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3757 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3758 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3759 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3760 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3761 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3762 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3763 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3764 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3765 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3766 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3767 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3768 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3769 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3770 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3771 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3772 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3773 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3774 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3775 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3776 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3777 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3778 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3779 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3780 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3781 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3782 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3783 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3784 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3785 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3786 AVDD|AVSS|VDD|VSS IREF \$19851 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3787 \$19851 IREF AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3788 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3789 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3790 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3791 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3792 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3793 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3794 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3795 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3796 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3797 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3798 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3799 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3800 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3801 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3802 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3803 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3804 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3805 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3806 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3807 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3808 AVDD|AVSS|VDD|VSS \$12262 \$19584 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3809 \$19584 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3810 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3811 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3812 AVDD|AVSS|VDD|VSS \$12262 \$19852 AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3813 \$19852 \$12262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS pfet_03v3 L=2U W=2U
+ AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3814 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3815 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3816 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3817 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3818 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3819 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3820 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3821 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3822 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3823 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3824 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3825 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3826 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3827 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3828 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3829 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3830 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3831 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3832 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3833 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3834 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3835 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3836 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3837 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3838 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3839 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3840 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3841 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3842 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3843 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3844 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3845 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3846 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3847 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3848 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3849 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3850 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3851 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3852 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3853 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3854 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3855 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3856 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3857 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3858 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3859 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3860 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3861 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3862 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3863 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3864 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3865 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3866 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS
+ pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3867 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3868 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3869 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3870 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3871 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3872 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3873 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3874 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3875 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3876 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3877 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3878 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3879 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3880 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3881 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3882 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3883 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3884 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3885 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3886 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3887 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3888 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3889 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3890 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3891 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3892 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3893 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3894 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3895 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3896 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3897 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3898 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3899 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3900 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3901 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3902 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3903 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3904 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3905 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3906 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3907 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3908 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3909 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3910 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3911 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3912 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3913 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3914 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3915 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3916 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3917 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3918 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3919 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3920 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3921 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3922 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3923 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3924 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3925 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3926 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3927 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3928 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3929 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3930 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3931 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3932 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3933 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3934 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3935 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3936 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3937 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3938 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3939 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3940 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3941 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3942 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3943 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3944 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3945 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3946 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3947 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3948 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3949 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3950 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3951 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3952 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3953 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3954 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3955 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3956 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3957 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3958 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3959 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3960 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3961 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3962 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3963 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3964 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3965 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3966 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3967 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3968 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3969 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3970 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3971 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3972 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3973 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3974 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3975 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3976 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3977 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3978 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3979 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3980 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3981 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3982 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3983 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3984 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3985 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3986 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3987 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3988 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3989 \$886 \$916 \$917 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$3990 \$866 \$916 \$886 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$3991 \$887 \$258 \$866 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$3992 \$172 \$258 \$887 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$3993 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3994 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3995 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3996 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3997 \$888 \$917 \$138 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$3998 \$258 \$917 \$888 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$3999 \$889 \$917 \$258 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4000 \$115 \$917 \$889 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4001 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4002 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4003 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4004 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4005 \$890 \$257 \$24 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4006 AVDD|AVSS|VDD|VSS \$257 \$890 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4007 \$891 \$257 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4008 \$257 \$257 \$891 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4009 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4010 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4011 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4012 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4013 \$892 \$918 \$919 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4014 \$867 \$918 \$892 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4015 \$893 \$260 \$867 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4016 \$174 \$260 \$893 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4017 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4018 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4019 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4020 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4021 \$894 \$919 \$146 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4022 \$260 \$919 \$894 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4023 \$895 \$919 \$260 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4024 \$116 \$919 \$895 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4025 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4026 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4027 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4028 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4029 \$896 \$259 \$25 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4030 AVDD|AVSS|VDD|VSS \$259 \$896 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4031 \$897 \$259 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4032 \$259 \$259 \$897 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4033 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4034 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4035 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4036 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4037 \$898 \$920 \$921 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4038 \$868 \$920 \$898 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4039 \$899 \$262 \$868 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4040 \$176 \$262 \$899 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4041 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4042 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4043 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4044 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4045 \$900 \$921 \$153 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4046 \$262 \$921 \$900 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4047 \$901 \$921 \$262 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4048 \$117 \$921 \$901 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4049 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4050 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4051 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4052 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4053 \$902 \$261 \$26 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4054 AVDD|AVSS|VDD|VSS \$261 \$902 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4055 \$903 \$261 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4056 \$261 \$261 \$903 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4057 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4058 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4059 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4060 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4061 \$904 \$922 \$923 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4062 \$869 \$922 \$904 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4063 \$905 \$264 \$869 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4064 \$178 \$264 \$905 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4065 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4066 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4067 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4068 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4069 \$906 \$923 \$160 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4070 \$264 \$923 \$906 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4071 \$907 \$923 \$264 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4072 \$118 \$923 \$907 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4073 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4074 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4075 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4076 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4077 \$908 \$263 \$27 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4078 AVDD|AVSS|VDD|VSS \$263 \$908 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4079 \$909 \$263 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4080 \$263 \$263 \$909 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4081 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4082 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4083 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4084 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4085 \$910 \$924 \$925 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4086 \$870 \$924 \$910 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4087 \$911 \$266 \$870 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4088 \$180 \$266 \$911 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4089 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4090 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4091 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4092 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4093 \$912 \$925 \$168 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4094 \$266 \$925 \$912 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4095 \$913 \$925 \$266 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4096 \$119 \$925 \$913 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4097 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4098 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4099 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4100 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4101 \$914 \$265 \$28 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4102 AVDD|AVSS|VDD|VSS \$265 \$914 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4103 \$915 \$265 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4104 \$265 \$265 \$915 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4105 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4106 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4107 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4108 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4109 \$1041 \$258 \$172 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4110 \$866 \$258 \$1041 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4111 \$1042 \$916 \$866 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4112 \$917 \$916 \$1042 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4113 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4114 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4115 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4116 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4117 \$1043 \$917 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4118 \$916 \$917 \$1043 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4119 \$1044 \$917 \$916 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4120 AVDD|AVSS|VDD|VSS \$917 \$1044 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4121 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4122 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4123 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4124 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4125 \$1045 \$257 \$257 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4126 AVDD|AVSS|VDD|VSS \$257 \$1045 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4127 \$1046 \$257 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4128 \$24 \$257 \$1046 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4129 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4130 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4131 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4132 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4133 \$1047 \$260 \$174 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4134 \$867 \$260 \$1047 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4135 \$1048 \$918 \$867 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4136 \$919 \$918 \$1048 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4137 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4138 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4139 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4140 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4141 \$1049 \$919 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4142 \$918 \$919 \$1049 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4143 \$1050 \$919 \$918 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4144 AVDD|AVSS|VDD|VSS \$919 \$1050 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4145 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4146 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4147 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4148 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4149 \$1051 \$259 \$259 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4150 AVDD|AVSS|VDD|VSS \$259 \$1051 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4151 \$1052 \$259 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4152 \$25 \$259 \$1052 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4153 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4154 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4155 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4156 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4157 \$1053 \$262 \$176 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4158 \$868 \$262 \$1053 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4159 \$1054 \$920 \$868 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4160 \$921 \$920 \$1054 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4161 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4162 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4163 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4164 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4165 \$1055 \$921 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4166 \$920 \$921 \$1055 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4167 \$1056 \$921 \$920 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4168 AVDD|AVSS|VDD|VSS \$921 \$1056 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4169 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4170 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4171 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4172 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4173 \$1057 \$261 \$261 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4174 AVDD|AVSS|VDD|VSS \$261 \$1057 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4175 \$1058 \$261 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4176 \$26 \$261 \$1058 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4177 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4178 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4179 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4180 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4181 \$1059 \$264 \$178 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4182 \$869 \$264 \$1059 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4183 \$1060 \$922 \$869 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4184 \$923 \$922 \$1060 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4185 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4186 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4187 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4188 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4189 \$1061 \$923 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4190 \$922 \$923 \$1061 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4191 \$1062 \$923 \$922 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4192 AVDD|AVSS|VDD|VSS \$923 \$1062 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4193 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4194 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4195 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4196 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4197 \$1063 \$263 \$263 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4198 AVDD|AVSS|VDD|VSS \$263 \$1063 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4199 \$1064 \$263 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4200 \$27 \$263 \$1064 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4201 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4202 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4203 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4204 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4205 \$1065 \$266 \$180 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4206 \$870 \$266 \$1065 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4207 \$1066 \$924 \$870 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4208 \$925 \$924 \$1066 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4209 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4210 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4211 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4212 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4213 \$1067 \$925 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4214 \$924 \$925 \$1067 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4215 \$1068 \$925 \$924 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4216 AVDD|AVSS|VDD|VSS \$925 \$1068 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4217 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4218 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4219 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4220 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4221 \$1069 \$265 \$265 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4222 AVDD|AVSS|VDD|VSS \$265 \$1069 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4223 \$1070 \$265 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4224 \$28 \$265 \$1070 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4225 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4226 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4227 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4228 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4229 \$1176 \$916 \$917 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4230 \$866 \$916 \$1176 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4231 \$1177 \$258 \$866 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4232 \$172 \$258 \$1177 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4233 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4234 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4235 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4236 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4237 \$1178 \$917 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4238 \$916 \$917 \$1178 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4239 \$1179 \$917 \$916 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4240 AVDD|AVSS|VDD|VSS \$917 \$1179 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4241 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4242 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4243 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4244 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4245 \$1180 \$257 \$24 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4246 AVDD|AVSS|VDD|VSS \$257 \$1180 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4247 \$1181 \$257 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4248 \$257 \$257 \$1181 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4249 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4250 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4251 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4252 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4253 \$1182 \$918 \$919 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4254 \$867 \$918 \$1182 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4255 \$1183 \$260 \$867 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4256 \$174 \$260 \$1183 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4257 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4258 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4259 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4260 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4261 \$1184 \$919 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4262 \$918 \$919 \$1184 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4263 \$1185 \$919 \$918 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4264 AVDD|AVSS|VDD|VSS \$919 \$1185 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4265 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4266 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4267 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4268 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4269 \$1186 \$259 \$25 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4270 AVDD|AVSS|VDD|VSS \$259 \$1186 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4271 \$1187 \$259 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4272 \$259 \$259 \$1187 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4273 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4274 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4275 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4276 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4277 \$1188 \$920 \$921 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4278 \$868 \$920 \$1188 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4279 \$1189 \$262 \$868 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4280 \$176 \$262 \$1189 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4281 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4282 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4283 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4284 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4285 \$1190 \$921 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4286 \$920 \$921 \$1190 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4287 \$1191 \$921 \$920 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4288 AVDD|AVSS|VDD|VSS \$921 \$1191 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4289 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4290 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4291 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4292 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4293 \$1192 \$261 \$26 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4294 AVDD|AVSS|VDD|VSS \$261 \$1192 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4295 \$1193 \$261 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4296 \$261 \$261 \$1193 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4297 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4298 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4299 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4300 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4301 \$1194 \$922 \$923 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4302 \$869 \$922 \$1194 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4303 \$1195 \$264 \$869 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4304 \$178 \$264 \$1195 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4305 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4306 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4307 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4308 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4309 \$1196 \$923 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4310 \$922 \$923 \$1196 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4311 \$1197 \$923 \$922 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4312 AVDD|AVSS|VDD|VSS \$923 \$1197 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4313 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4314 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4315 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4316 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4317 \$1198 \$263 \$27 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4318 AVDD|AVSS|VDD|VSS \$263 \$1198 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4319 \$1199 \$263 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4320 \$263 \$263 \$1199 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4321 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4322 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4323 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4324 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4325 \$1200 \$924 \$925 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4326 \$870 \$924 \$1200 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4327 \$1201 \$266 \$870 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4328 \$180 \$266 \$1201 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4329 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4330 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4331 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4332 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4333 \$1202 \$925 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4334 \$924 \$925 \$1202 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4335 \$1203 \$925 \$924 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4336 AVDD|AVSS|VDD|VSS \$925 \$1203 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4337 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4338 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4339 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4340 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4341 \$1204 \$265 \$28 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4342 AVDD|AVSS|VDD|VSS \$265 \$1204 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4343 \$1205 \$265 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4344 \$265 \$265 \$1205 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4345 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4346 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4347 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4348 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4349 \$1321 \$258 \$172 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4350 \$866 \$258 \$1321 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4351 \$1322 \$916 \$866 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4352 \$917 \$916 \$1322 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4353 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4354 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4355 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4356 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4357 \$1323 \$917 \$115 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4358 \$258 \$917 \$1323 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4359 \$1324 \$917 \$258 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4360 \$138 \$917 \$1324 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4361 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4362 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4363 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4364 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4365 \$1325 \$257 \$257 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4366 AVDD|AVSS|VDD|VSS \$257 \$1325 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4367 \$1326 \$257 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4368 \$24 \$257 \$1326 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4369 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4370 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4371 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4372 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4373 \$1327 \$260 \$174 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4374 \$867 \$260 \$1327 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4375 \$1328 \$918 \$867 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4376 \$919 \$918 \$1328 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4377 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4378 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4379 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4380 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4381 \$1329 \$919 \$116 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4382 \$260 \$919 \$1329 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4383 \$1330 \$919 \$260 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4384 \$146 \$919 \$1330 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4385 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4386 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4387 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4388 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4389 \$1331 \$259 \$259 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4390 AVDD|AVSS|VDD|VSS \$259 \$1331 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4391 \$1332 \$259 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4392 \$25 \$259 \$1332 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4393 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4394 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4395 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4396 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4397 \$1333 \$262 \$176 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4398 \$868 \$262 \$1333 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4399 \$1334 \$920 \$868 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4400 \$921 \$920 \$1334 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4401 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4402 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4403 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4404 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4405 \$1335 \$921 \$117 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4406 \$262 \$921 \$1335 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4407 \$1336 \$921 \$262 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4408 \$153 \$921 \$1336 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4409 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4410 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4411 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4412 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4413 \$1337 \$261 \$261 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4414 AVDD|AVSS|VDD|VSS \$261 \$1337 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4415 \$1338 \$261 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4416 \$26 \$261 \$1338 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4417 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4418 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4419 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4420 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4421 \$1339 \$264 \$178 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4422 \$869 \$264 \$1339 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4423 \$1340 \$922 \$869 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4424 \$923 \$922 \$1340 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4425 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4426 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4427 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4428 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4429 \$1341 \$923 \$118 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4430 \$264 \$923 \$1341 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4431 \$1342 \$923 \$264 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4432 \$160 \$923 \$1342 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4433 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4434 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4435 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4436 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4437 \$1343 \$263 \$263 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4438 AVDD|AVSS|VDD|VSS \$263 \$1343 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4439 \$1344 \$263 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4440 \$27 \$263 \$1344 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4441 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4442 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4443 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4444 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4445 \$1345 \$266 \$180 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4446 \$870 \$266 \$1345 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4447 \$1346 \$924 \$870 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4448 \$925 \$924 \$1346 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4449 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4450 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4451 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4452 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4453 \$1347 \$925 \$119 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4454 \$266 \$925 \$1347 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4455 \$1348 \$925 \$266 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4456 \$168 \$925 \$1348 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4457 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4458 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4459 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4460 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4461 \$1349 \$265 \$265 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4462 AVDD|AVSS|VDD|VSS \$265 \$1349 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4463 \$1350 \$265 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$4464 \$28 \$265 \$1350 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4465 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4466 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4467 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4468 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4469 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4470 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4471 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4472 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4473 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4474 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4475 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4476 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4477 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4478 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4479 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4480 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4481 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4482 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4483 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4484 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4485 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4486 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4487 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4488 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4489 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4490 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4491 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4492 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4493 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4494 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4495 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4496 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4497 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4498 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4499 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4500 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4501 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4502 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4503 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4504 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4505 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4506 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4507 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4508 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4509 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4510 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4511 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4512 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4513 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4514 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4515 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4516 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4517 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4518 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4519 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4520 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4521 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4522 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4523 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4524 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4525 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4526 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4527 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4528 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4529 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4530 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4531 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4532 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4533 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4534 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4535 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4536 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4537 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4538 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4539 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4540 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4541 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4542 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4543 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4544 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4545 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4546 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4547 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4548 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4549 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4550 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4551 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4552 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4553 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4554 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4555 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4556 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4557 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4558 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4559 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4560 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4561 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4562 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4563 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4564 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4565 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4566 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4567 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4568 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4569 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4570 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4571 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4572 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4575 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4576 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4577 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4578 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4579 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4580 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4581 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4582 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4583 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4584 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4585 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4586 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4587 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4588 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4589 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4590 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4591 \$1782 \$1774 \$1781 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4592 \$916 \$1774 \$1782 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4593 \$1784 \$1774 \$1783 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4594 \$1785 \$1774 \$1784 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4595 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4596 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4597 \$1786 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4598 \$1787 \$1774 \$1786 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4599 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4600 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4601 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4602 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4603 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4604 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4605 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4606 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4607 \$1789 \$1774 \$1788 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4608 \$918 \$1774 \$1789 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4609 \$1791 \$1774 \$1790 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4610 \$1792 \$1774 \$1791 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4611 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4612 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4613 \$1793 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4614 \$1794 \$1774 \$1793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4615 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4616 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4617 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4618 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4619 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4620 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4621 \$1796 \$1774 \$1795 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4622 \$920 \$1774 \$1796 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4623 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4624 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4625 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4626 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4627 \$1798 \$1774 \$1797 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4628 \$1799 \$1774 \$1798 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4629 \$1800 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4630 \$1801 \$1774 \$1800 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4631 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4632 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4633 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4634 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4635 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4636 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4637 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4638 \$1958 \$1731 \$1802 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4639 \$1959 \$1731 \$1958 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4640 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4641 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4642 \$1803 \$1731 \$1802 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4643 \$1732 \$1731 \$1803 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4644 \$1961 \$1731 \$1960 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4645 \$1805 \$1731 \$1961 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4646 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4647 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4648 \$1804 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4649 \$1805 \$1731 \$1804 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4650 \$1963 \$1731 \$1962 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4651 \$1807 \$1731 \$1963 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4652 \$1806 \$1731 \$1732 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4653 \$1807 \$1731 \$1806 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4654 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4655 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4656 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4657 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4658 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4659 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4660 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4661 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4662 \$1964 \$1731 \$1808 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4663 \$1965 \$1731 \$1964 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4664 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4665 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4666 \$1809 \$1731 \$1808 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4667 \$1733 \$1731 \$1809 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4668 \$1810 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4669 \$1811 \$1731 \$1810 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4670 \$1967 \$1731 \$1966 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4671 \$1811 \$1731 \$1967 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4672 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4673 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4674 \$1969 \$1731 \$1968 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4675 \$1813 \$1731 \$1969 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4676 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4677 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4678 \$1812 \$1731 \$1733 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4679 \$1813 \$1731 \$1812 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4680 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4681 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4682 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4683 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4684 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4685 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4686 \$1815 \$1731 \$1814 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4687 \$1734 \$1731 \$1815 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4688 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4689 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4690 \$1970 \$1731 \$1814 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4691 \$1971 \$1731 \$1970 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4692 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4693 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4694 \$1973 \$1731 \$1972 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4695 \$1817 \$1731 \$1973 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4696 \$1816 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4697 \$1817 \$1731 \$1816 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4698 \$1818 \$1731 \$1734 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4699 \$1819 \$1731 \$1818 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4700 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4701 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4702 \$1975 \$1731 \$1974 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4703 \$1819 \$1731 \$1975 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4704 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4705 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4706 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4707 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4708 \$1940 \$1774 \$1781 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4709 \$1941 \$1774 \$1940 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4710 \$1943 \$1774 \$1942 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4711 \$1785 \$1774 \$1943 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4712 \$1945 \$1774 \$1944 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4713 \$1787 \$1774 \$1945 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4714 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4715 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4716 \$1946 \$1774 \$1788 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4717 \$1947 \$1774 \$1946 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4718 \$1949 \$1774 \$1948 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4719 \$1792 \$1774 \$1949 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4720 \$1951 \$1774 \$1950 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4721 \$1794 \$1774 \$1951 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4722 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4723 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4724 \$1952 \$1774 \$1795 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4725 \$1953 \$1774 \$1952 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4726 \$1955 \$1774 \$1954 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4727 \$1799 \$1774 \$1955 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4728 \$1957 \$1774 \$1956 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4729 \$1801 \$1774 \$1957 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4730 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4731 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4732 \$2130 \$1774 \$2129 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4733 \$1941 \$1774 \$2130 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4734 \$2131 \$1774 \$1942 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4735 \$2132 \$1774 \$2131 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4736 \$2133 \$1774 \$1944 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4737 \$2134 \$1774 \$2133 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4738 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4739 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4740 \$2136 \$1774 \$2135 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4741 \$1947 \$1774 \$2136 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4742 \$2137 \$1774 \$1948 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4743 \$2138 \$1774 \$2137 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4744 \$2139 \$1774 \$1950 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4745 \$2140 \$1774 \$2139 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4746 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4747 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4748 \$2142 \$1774 \$2141 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4749 \$1953 \$1774 \$2142 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4750 \$2143 \$1774 \$1954 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4751 \$2144 \$1774 \$2143 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4752 \$2145 \$1774 \$1956 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4753 \$2146 \$1774 \$2145 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4754 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4755 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4756 \$2103 \$1731 \$2102 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4757 \$1959 \$1731 \$2103 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4758 \$2104 \$1731 \$1960 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4759 \$2048 \$1731 \$2104 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4760 \$2105 \$1731 \$1962 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4761 \$2106 \$1731 \$2105 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4762 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4763 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4764 \$2108 \$1731 \$2107 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4765 \$1965 \$1731 \$2108 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4766 \$2109 \$1731 \$1966 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4767 \$2049 \$1731 \$2109 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4768 \$2110 \$1731 \$1968 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4769 \$2111 \$1731 \$2110 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4770 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4771 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4772 \$2113 \$1731 \$2112 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4773 \$1971 \$1731 \$2113 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4774 \$2114 \$1731 \$1972 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4775 \$2050 \$1731 \$2114 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4776 \$2115 \$1731 \$1974 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4777 \$2116 \$1731 \$2115 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4778 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4779 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4780 \$2266 \$1774 \$2129 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4781 \$2267 \$1774 \$2266 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4782 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4783 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4784 \$2269 \$1774 \$2268 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4785 \$2134 \$1774 \$2269 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4786 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4787 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4788 \$2270 \$1774 \$2135 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4789 \$2271 \$1774 \$2270 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4790 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4791 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4792 \$2273 \$1774 \$2272 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4793 \$2140 \$1774 \$2273 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4794 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4795 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4796 \$2274 \$1774 \$2141 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4797 \$2275 \$1774 \$2274 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4798 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4799 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4800 \$2277 \$1774 \$2276 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4801 \$2146 \$1774 \$2277 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4802 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4803 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4804 \$2278 \$1731 \$2102 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4805 \$2279 \$1731 \$2278 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4806 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4807 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4808 \$2281 \$1731 \$2280 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4809 \$2106 \$1731 \$2281 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4810 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4811 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4812 \$2282 \$1731 \$2107 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4813 \$2283 \$1731 \$2282 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4814 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4815 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4816 \$2285 \$1731 \$2284 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4817 \$2111 \$1731 \$2285 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4818 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4819 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4820 \$2286 \$1731 \$2112 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4821 \$2287 \$1731 \$2286 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4822 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4823 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4824 \$2289 \$1731 \$2288 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4825 \$2116 \$1731 \$2289 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4826 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4827 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4828 \$2407 \$1774 \$866 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4829 \$1783 \$1774 \$2407 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4830 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4831 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4832 \$2408 \$1774 \$2132 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4833 \$2409 \$1774 \$2408 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4834 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4835 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4836 \$2410 \$1774 \$867 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4837 \$1790 \$1774 \$2410 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4838 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4839 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4840 \$2411 \$1774 \$2138 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4841 \$2412 \$1774 \$2411 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4842 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4843 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4844 \$2413 \$1774 \$868 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4845 \$1797 \$1774 \$2413 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4846 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4847 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4848 \$2414 \$1774 \$2144 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4849 \$2415 \$1774 \$2414 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4850 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4851 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4852 \$2416 \$1731 \$5350 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4853 \$2417 \$1731 \$2416 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4854 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4855 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4856 \$2418 \$1731 \$2443 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4857 \$2048 \$1731 \$2418 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4858 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4859 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4860 \$2419 \$1731 \$5351 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4861 \$2420 \$1731 \$2419 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4862 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4863 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4864 \$2421 \$1731 \$2444 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4865 \$2049 \$1731 \$2421 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4866 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4867 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4868 \$2422 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4869 \$2423 \$1731 \$2422 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4870 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4871 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4872 \$2424 \$1731 \$2445 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4873 \$2050 \$1731 \$2424 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4874 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4875 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4876 \$2637 \$1774 \$2636 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4877 \$2267 \$1774 \$2637 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4878 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4879 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4880 \$2638 \$1774 \$2268 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4881 \$2639 \$1774 \$2638 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4882 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4883 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4884 \$2641 \$1774 \$2640 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4885 \$2271 \$1774 \$2641 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4886 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4887 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4888 \$2642 \$1774 \$2272 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4889 \$2643 \$1774 \$2642 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4890 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4891 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4892 \$2645 \$1774 \$2644 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4893 \$2275 \$1774 \$2645 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4894 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4895 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4896 \$2646 \$1774 \$2276 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4897 \$2647 \$1774 \$2646 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4898 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4899 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4900 \$2589 \$1731 \$2588 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4901 \$2279 \$1731 \$2589 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4902 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4903 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4904 \$2590 \$1731 \$2280 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4905 \$2591 \$1731 \$2590 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4906 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4907 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4908 \$2593 \$1731 \$2592 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4909 \$2283 \$1731 \$2593 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4910 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4911 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4912 \$2594 \$1731 \$2284 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4913 \$2595 \$1731 \$2594 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4914 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4915 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4916 \$2597 \$1731 \$2596 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4917 \$2287 \$1731 \$2597 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4918 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4919 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$4920 \$2598 \$1731 \$2288 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4921 \$2599 \$1731 \$2598 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4922 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4923 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4924 \$2906 \$1774 \$2636 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4925 \$2907 \$1774 \$2906 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4926 \$2909 \$1774 \$2908 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4927 \$2409 \$1774 \$2909 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4928 \$2911 \$1774 \$2910 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4929 \$2639 \$1774 \$2911 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4930 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4931 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4932 \$2912 \$1774 \$2640 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4933 \$2913 \$1774 \$2912 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4934 \$2915 \$1774 \$2914 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4935 \$2412 \$1774 \$2915 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4936 \$2917 \$1774 \$2916 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4937 \$2643 \$1774 \$2917 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4938 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4939 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4940 \$2918 \$1774 \$2644 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4941 \$2919 \$1774 \$2918 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4942 \$2921 \$1774 \$2920 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4943 \$2415 \$1774 \$2921 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4944 \$2923 \$1774 \$2922 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4945 \$2647 \$1774 \$2923 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4946 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4947 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4948 \$2924 \$1731 \$2588 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4949 \$2925 \$1731 \$2924 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4950 \$2927 \$1731 \$2926 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4951 \$2443 \$1731 \$2927 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4952 \$2929 \$1731 \$2928 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4953 \$2591 \$1731 \$2929 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4954 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4955 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4956 \$2930 \$1731 \$2592 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4957 \$2931 \$1731 \$2930 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4958 \$2933 \$1731 \$2932 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4959 \$2444 \$1731 \$2933 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4960 \$2935 \$1731 \$2934 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4961 \$2595 \$1731 \$2935 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4962 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4963 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4964 \$2936 \$1731 \$2596 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4965 \$2937 \$1731 \$2936 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4966 \$2939 \$1731 \$2938 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4967 \$2445 \$1731 \$2939 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4968 \$2941 \$1731 \$2940 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4969 \$2599 \$1731 \$2941 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4970 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4971 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4972 \$3172 \$1774 \$3171 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4973 \$2907 \$1774 \$3172 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4974 \$3173 \$1774 \$2908 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4975 \$3174 \$1774 \$3173 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4976 \$3175 \$1774 \$2910 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4977 \$3176 \$1774 \$3175 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4978 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4979 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4980 \$3178 \$1774 \$3177 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4981 \$2913 \$1774 \$3178 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4982 \$3179 \$1774 \$2914 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4983 \$3180 \$1774 \$3179 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4984 \$3181 \$1774 \$2916 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4985 \$3182 \$1774 \$3181 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4986 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4987 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4988 \$3184 \$1774 \$3183 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4989 \$2919 \$1774 \$3184 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4990 \$3185 \$1774 \$2920 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4991 \$3186 \$1774 \$3185 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4992 \$3187 \$1774 \$2922 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4993 \$3188 \$1774 \$3187 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4994 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4995 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4996 \$3190 \$1731 \$3189 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4997 \$2925 \$1731 \$3190 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$4998 \$3191 \$1731 \$2926 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$4999 \$3192 \$1731 \$3191 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5000 \$3193 \$1731 \$2928 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5001 \$3194 \$1731 \$3193 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5002 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5003 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5004 \$3196 \$1731 \$3195 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5005 \$2931 \$1731 \$3196 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5006 \$3197 \$1731 \$2932 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5007 \$3198 \$1731 \$3197 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5008 \$3199 \$1731 \$2934 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5009 \$3200 \$1731 \$3199 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5010 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5011 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5012 \$3202 \$1731 \$3201 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5013 \$2937 \$1731 \$3202 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5014 \$3203 \$1731 \$2938 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5015 \$3204 \$1731 \$3203 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5016 \$3205 \$1731 \$2940 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5017 \$3206 \$1731 \$3205 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5018 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5019 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5020 \$3360 \$1774 \$3171 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5021 \$3361 \$1774 \$3360 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5022 \$3362 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5023 \$3174 \$1774 \$3362 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5024 \$3363 \$1774 \$3361 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5025 \$3176 \$1774 \$3363 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5026 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5027 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5028 \$3364 \$1774 \$3177 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5029 \$3365 \$1774 \$3364 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5030 \$3366 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5031 \$3180 \$1774 \$3366 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5032 \$3367 \$1774 \$3365 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5033 \$3182 \$1774 \$3367 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5034 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5035 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5036 \$3368 \$1774 \$3183 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5037 \$3369 \$1774 \$3368 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5038 \$3370 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5039 \$3186 \$1774 \$3370 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5040 \$3371 \$1774 \$3369 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5041 \$3188 \$1774 \$3371 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5042 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5043 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5044 \$3345 \$1731 \$3189 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5045 \$3346 \$1731 \$3345 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5046 \$3347 \$1731 \$2417 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5047 \$3192 \$1731 \$3347 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5048 \$3348 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5049 \$3194 \$1731 \$3348 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5050 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5051 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5052 \$3349 \$1731 \$3195 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5053 \$3350 \$1731 \$3349 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5054 \$3351 \$1731 \$2420 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5055 \$3198 \$1731 \$3351 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5056 \$3352 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5057 \$3200 \$1731 \$3352 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5058 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5059 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5060 \$3353 \$1731 \$3201 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5061 CMOUTN \$1731 \$3353 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5062 \$3355 \$1731 \$2423 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5063 \$3204 \$1731 \$3355 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5064 \$3356 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5065 \$3206 \$1731 \$3356 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5066 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5067 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5068 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5069 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5070 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5071 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5072 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5073 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5074 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5075 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5076 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5077 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5078 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5079 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5080 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5081 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5082 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5083 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5084 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5085 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5086 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5087 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5088 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5089 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5090 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5091 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5092 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5093 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5094 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5095 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5096 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5097 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5098 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5099 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5100 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5101 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5102 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5103 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5104 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5105 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5106 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5107 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5108 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5109 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5110 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5111 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5112 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5113 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5114 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5115 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5116 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5117 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5118 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5119 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5120 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5121 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5122 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5123 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5124 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5125 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5126 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5127 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5128 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5129 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5130 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5131 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5132 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5133 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5134 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5135 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5136 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5137 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5138 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5139 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5140 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5141 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5142 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5143 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5144 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5145 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5146 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5147 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5148 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5149 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5150 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5151 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5152 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5153 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5154 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5155 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5156 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5157 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5158 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5159 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5160 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5161 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5162 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5163 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5164 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5165 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5166 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5167 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5168 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5169 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5170 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5171 \$3462 ISBCS ISBCS gf180mcu_gnd nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5172 AVDD|AVSS|VDD|VSS ISBCS \$3462 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5173 \$3549 ISBCS \$1573 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5174 AVDD|AVSS|VDD|VSS ISBCS \$3549 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5175 \$3463 ISBCS AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=6U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$5176 \$1574 ISBCS \$3463 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5177 \$3550 ISBCS AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=6U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$5178 \$4383 ISBCS \$3550 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5179 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5180 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5181 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5182 \$3699 \$1774 \$3698 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5183 \$922 \$1774 \$3699 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5184 \$3701 \$1774 \$3700 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5185 \$3702 \$1774 \$3701 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5186 \$3703 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5187 \$3704 \$1774 \$3703 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5188 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5189 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5190 \$3706 \$1774 \$3705 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5191 \$924 \$1774 \$3706 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5192 \$3708 \$1774 \$3707 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5193 \$3709 \$1774 \$3708 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5194 \$3710 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5195 \$3711 \$1774 \$3710 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5196 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5197 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5198 \$3713 \$1774 \$3712 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5199 AVDD|AVSS|VDD|VSS \$1774 \$3713 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5200 \$3715 \$1774 \$3714 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5201 \$3716 \$1774 \$3715 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5202 \$3717 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5203 \$3718 \$1774 \$3717 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5204 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5205 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5206 \$3720 \$1731 \$3719 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5207 \$3673 \$1731 \$3720 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5208 \$3721 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5209 \$3722 \$1731 \$3721 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5210 \$3723 \$1731 \$3673 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5211 \$3724 \$1731 \$3723 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5212 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5213 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5214 \$3726 \$1731 \$3725 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5215 \$3674 \$1731 \$3726 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5216 \$3727 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5217 \$3728 \$1731 \$3727 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5218 \$3729 \$1731 \$3674 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5219 \$3730 \$1731 \$3729 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5220 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5221 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5222 \$3732 \$1731 \$3731 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5223 \$3675 \$1731 \$3732 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5224 \$3733 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5225 \$3734 \$1731 \$3733 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5226 \$3735 \$1731 \$3675 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5227 \$3736 \$1731 \$3735 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5228 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5229 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5230 \$3629 ISBCS \$1573 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5231 AVDD|AVSS|VDD|VSS ISBCS \$3629 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5232 \$3630 ISBCS AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=6U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$5233 \$4383 ISBCS \$3630 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5234 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5235 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5236 \$3862 \$1774 \$3698 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5237 \$3863 \$1774 \$3862 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5238 \$3865 \$1774 \$3864 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5239 \$3702 \$1774 \$3865 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5240 \$3867 \$1774 \$3866 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5241 \$3704 \$1774 \$3867 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5242 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5243 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5244 \$3868 \$1774 \$3705 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5245 \$3869 \$1774 \$3868 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5246 \$3871 \$1774 \$3870 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5247 \$3709 \$1774 \$3871 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5248 \$3873 \$1774 \$3872 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5249 \$3711 \$1774 \$3873 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5250 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5251 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5252 \$3874 \$1774 \$3712 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5253 \$3875 \$1774 \$3874 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5254 \$3877 \$1774 \$3876 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5255 \$3716 \$1774 \$3877 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5256 \$3879 \$1774 \$3878 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5257 \$3718 \$1774 \$3879 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5258 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5259 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5260 \$3880 \$1731 \$3719 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5261 \$3881 \$1731 \$3880 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5262 \$3883 \$1731 \$3882 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5263 \$3722 \$1731 \$3883 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5264 \$3885 \$1731 \$3884 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5265 \$3724 \$1731 \$3885 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5266 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5267 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5268 \$3886 \$1731 \$3725 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5269 \$3887 \$1731 \$3886 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5270 \$3889 \$1731 \$3888 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5271 \$3728 \$1731 \$3889 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5272 \$3891 \$1731 \$3890 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5273 \$3730 \$1731 \$3891 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5274 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5275 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5276 \$3892 \$1731 \$3731 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5277 \$3893 \$1731 \$3892 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5278 \$3895 \$1731 \$3894 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5279 \$3734 \$1731 \$3895 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5280 \$3897 \$1731 \$3896 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5281 \$3736 \$1731 \$3897 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5282 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5283 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5284 \$3811 ISBCS \$1574 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5285 AVDD|AVSS|VDD|VSS ISBCS \$3811 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5286 \$3812 ISBCS AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=6U W=2U AS=1.22P
+ AD=0.8P PS=5.22U PD=2.8U
M$5287 ISBCS ISBCS \$3812 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5288 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5289 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5290 \$4026 \$1774 \$4025 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5291 \$3863 \$1774 \$4026 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5292 \$4027 \$1774 \$3864 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5293 \$4028 \$1774 \$4027 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5294 \$4029 \$1774 \$3866 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5295 \$4030 \$1774 \$4029 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5296 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5297 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5298 \$4032 \$1774 \$4031 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5299 \$3869 \$1774 \$4032 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5300 \$4033 \$1774 \$3870 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5301 \$4034 \$1774 \$4033 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5302 \$4035 \$1774 \$3872 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5303 \$4036 \$1774 \$4035 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5304 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5305 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5306 \$4038 \$1774 \$4037 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5307 \$3875 \$1774 \$4038 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5308 \$4039 \$1774 \$3876 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5309 \$4040 \$1774 \$4039 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5310 \$4041 \$1774 \$3878 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5311 \$4042 \$1774 \$4041 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5312 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5313 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5314 \$4044 \$1731 \$4043 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5315 \$3881 \$1731 \$4044 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5316 \$4045 \$1731 \$3882 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5317 \$4006 \$1731 \$4045 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5318 \$4046 \$1731 \$3884 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5319 \$4047 \$1731 \$4046 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5320 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5321 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5322 \$4049 \$1731 \$4048 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5323 \$3887 \$1731 \$4049 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5324 \$4050 \$1731 \$3888 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5325 \$4007 \$1731 \$4050 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5326 \$4051 \$1731 \$3890 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5327 \$4052 \$1731 \$4051 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5328 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5329 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5330 \$4054 \$1731 \$4053 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5331 \$3893 \$1731 \$4054 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5332 \$4055 \$1731 \$3894 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5333 \$4008 \$1731 \$4055 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5334 \$4056 \$1731 \$3896 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5335 \$4057 \$1731 \$4056 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5336 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5337 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5338 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5339 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5340 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5341 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5342 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5343 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5344 \$4198 \$1774 \$4025 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5345 \$4199 \$1774 \$4198 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5346 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5347 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5348 \$4201 \$1774 \$4200 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5349 \$4030 \$1774 \$4201 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5350 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5351 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5352 \$4202 \$1774 \$4031 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5353 \$4203 \$1774 \$4202 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5354 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5355 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5356 \$4205 \$1774 \$4204 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5357 \$4036 \$1774 \$4205 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5358 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5359 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5360 \$4206 \$1774 \$4037 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5361 \$4207 \$1774 \$4206 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5362 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5363 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5364 \$4209 \$1774 \$4208 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5365 \$4042 \$1774 \$4209 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5366 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5367 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5368 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5369 \$4371 \$1731 \$5347 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5370 \$4372 \$1731 \$4371 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5371 \$4210 \$1731 \$4043 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5372 \$4211 \$1731 \$4210 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5373 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5374 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5375 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5376 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5377 \$4213 \$1731 \$4212 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5378 \$4047 \$1731 \$4213 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5379 \$4373 \$1731 \$4380 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5380 \$4006 \$1731 \$4373 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5381 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5382 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5383 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5384 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5385 \$4374 \$1731 \$5348 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5386 \$4375 \$1731 \$4374 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5387 \$4214 \$1731 \$4048 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5388 \$4215 \$1731 \$4214 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5389 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5390 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5391 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5392 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5393 \$4217 \$1731 \$4216 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5394 \$4052 \$1731 \$4217 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5395 \$4376 \$1731 \$4381 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5396 \$4007 \$1731 \$4376 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5397 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5398 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5399 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5400 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5401 \$4377 \$1731 \$5349 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5402 \$4378 \$1731 \$4377 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5403 \$4218 \$1731 \$4053 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5404 \$4219 \$1731 \$4218 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5405 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5406 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5407 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5408 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5409 \$4221 \$1731 \$4220 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5410 \$4057 \$1731 \$4221 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5411 \$4379 \$1731 \$4382 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5412 \$4008 \$1731 \$4379 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5413 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5414 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5415 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5416 \$4362 \$1774 \$869 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5417 \$3700 \$1774 \$4362 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5418 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5419 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5420 \$4363 \$1774 \$4028 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5421 \$4364 \$1774 \$4363 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5422 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5423 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5424 \$4365 \$1774 \$870 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5425 \$3707 \$1774 \$4365 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5426 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5427 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5428 \$4366 \$1774 \$4034 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5429 \$4367 \$1774 \$4366 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5430 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5431 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5432 \$4368 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5433 \$3714 \$1774 \$4368 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5434 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5435 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5436 \$4369 \$1774 \$4040 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5437 \$4370 \$1774 \$4369 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5438 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5439 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5440 \$4522 \$1774 \$4521 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5441 \$4199 \$1774 \$4522 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5442 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5443 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5444 \$4523 \$1774 \$4200 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5445 \$4524 \$1774 \$4523 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5446 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5447 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5448 \$4526 \$1774 \$4525 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5449 \$4203 \$1774 \$4526 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5450 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5451 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5452 \$4527 \$1774 \$4204 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5453 \$4528 \$1774 \$4527 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5454 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5455 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5456 \$4530 \$1774 \$4529 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5457 \$4207 \$1774 \$4530 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5458 AVDD|AVSS|VDD|VSS \$1774 \$1774 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5459 \$1774 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5460 \$4531 \$1774 \$4208 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5461 \$4532 \$1774 \$4531 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5462 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5463 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5464 \$4534 \$1731 \$4533 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5465 \$4211 \$1731 \$4534 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5466 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5467 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5468 \$4535 \$1731 \$4212 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5469 \$4536 \$1731 \$4535 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5470 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5471 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5472 \$4538 \$1731 \$4537 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5473 \$4215 \$1731 \$4538 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5474 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5475 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5476 \$4539 \$1731 \$4216 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5477 \$4540 \$1731 \$4539 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5478 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5479 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5480 \$4542 \$1731 \$4541 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5481 \$4219 \$1731 \$4542 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5482 AVDD|AVSS|VDD|VSS \$1731 \$1731 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5483 \$1731 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5484 \$4543 \$1731 \$4220 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5485 \$4544 \$1731 \$4543 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5486 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5487 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5488 \$4694 \$1774 \$4521 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5489 \$4695 \$1774 \$4694 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5490 \$4697 \$1774 \$4696 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5491 \$4364 \$1774 \$4697 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5492 \$4699 \$1774 \$4698 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5493 \$4524 \$1774 \$4699 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5494 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5495 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5496 \$4700 \$1774 \$4525 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5497 \$4701 \$1774 \$4700 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5498 \$4703 \$1774 \$4702 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5499 \$4367 \$1774 \$4703 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5500 \$4705 \$1774 \$4704 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5501 \$4528 \$1774 \$4705 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5502 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5503 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5504 \$4706 \$1774 \$4529 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5505 \$4707 \$1774 \$4706 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5506 \$4709 \$1774 \$4708 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5507 \$4370 \$1774 \$4709 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5508 \$4711 \$1774 \$4710 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5509 \$4532 \$1774 \$4711 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5510 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5511 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5512 \$4712 \$1731 \$4533 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5513 \$4713 \$1731 \$4712 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5514 \$4715 \$1731 \$4714 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5515 \$4380 \$1731 \$4715 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5516 \$4717 \$1731 \$4716 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5517 \$4536 \$1731 \$4717 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5518 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5519 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5520 \$4718 \$1731 \$4537 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5521 \$4719 \$1731 \$4718 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5522 \$4721 \$1731 \$4720 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5523 \$4381 \$1731 \$4721 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5524 \$4723 \$1731 \$4722 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5525 \$4540 \$1731 \$4723 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5526 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5527 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5528 \$4724 \$1731 \$4541 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5529 \$4725 \$1731 \$4724 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5530 \$4727 \$1731 \$4726 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5531 \$4382 \$1731 \$4727 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5532 \$4729 \$1731 \$4728 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5533 \$4544 \$1731 \$4729 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5534 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5535 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5536 \$4870 \$1774 \$4869 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5537 \$4695 \$1774 \$4870 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5538 \$4871 \$1774 \$4696 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5539 \$4872 \$1774 \$4871 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5540 \$4873 \$1774 \$4698 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5541 \$4874 \$1774 \$4873 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5542 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5543 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5544 \$4876 \$1774 \$4875 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5545 \$4701 \$1774 \$4876 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5546 \$4877 \$1774 \$4702 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5547 \$4878 \$1774 \$4877 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5548 \$4879 \$1774 \$4704 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5549 \$4880 \$1774 \$4879 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5550 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5551 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5552 \$4882 \$1774 \$4881 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5553 \$4707 \$1774 \$4882 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5554 \$4883 \$1774 \$4708 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5555 \$4884 \$1774 \$4883 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5556 \$4885 \$1774 \$4710 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5557 \$4886 \$1774 \$4885 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5558 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5559 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5560 \$4888 \$1731 \$4887 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5561 \$4713 \$1731 \$4888 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5562 \$4889 \$1731 \$4714 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5563 \$4890 \$1731 \$4889 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5564 \$4891 \$1731 \$4716 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5565 \$4892 \$1731 \$4891 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5566 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5567 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5568 \$4894 \$1731 \$4893 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5569 \$4719 \$1731 \$4894 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5570 \$4895 \$1731 \$4720 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5571 \$4896 \$1731 \$4895 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5572 \$4897 \$1731 \$4722 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5573 \$4898 \$1731 \$4897 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5575 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5576 \$4900 \$1731 \$4899 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5577 \$4725 \$1731 \$4900 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5578 \$4901 \$1731 \$4726 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5579 \$4902 \$1731 \$4901 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5580 \$4903 \$1731 \$4728 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5581 \$4904 \$1731 \$4903 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5582 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5583 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5584 \$5010 \$1774 \$4869 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5585 \$5011 \$1774 \$5010 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5586 \$5012 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5587 \$4872 \$1774 \$5012 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5588 \$5013 \$1774 \$5011 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5589 \$4874 \$1774 \$5013 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5590 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5591 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5592 \$5014 \$1774 \$4875 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5593 \$5015 \$1774 \$5014 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5594 \$5016 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5595 \$4878 \$1774 \$5016 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5596 \$5017 \$1774 \$5015 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5597 \$4880 \$1774 \$5017 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5598 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5599 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5600 \$5018 \$1774 \$4881 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5601 \$5019 \$1774 \$5018 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5602 \$5020 \$1774 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5603 \$4884 \$1774 \$5020 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5604 \$5021 \$1774 \$5019 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5605 \$4886 \$1774 \$5021 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5606 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5607 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5608 \$5022 \$1731 \$4887 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5609 \$5023 \$1731 \$5022 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5610 \$5024 \$1731 \$4372 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5611 \$4890 \$1731 \$5024 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5612 \$5025 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5613 \$4892 \$1731 \$5025 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5614 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5615 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5616 \$5026 \$1731 \$4893 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5617 \$5027 \$1731 \$5026 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5618 \$5028 \$1731 \$4375 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5619 \$4896 \$1731 \$5028 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5620 \$5029 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5621 \$4898 \$1731 \$5029 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5622 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5623 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5624 \$5030 \$1731 \$4899 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5625 \$5031 \$1731 \$5030 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5626 \$5032 \$1731 \$4378 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5627 \$4902 \$1731 \$5032 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5628 \$5033 \$1731 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5629 \$4904 \$1731 \$5033 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5630 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5631 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5632 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5633 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5634 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5635 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5636 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5637 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5638 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5639 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5640 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5641 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5642 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5643 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5644 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5645 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5646 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5647 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5648 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5649 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5650 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5651 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5652 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5653 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5654 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5655 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5656 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5657 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5658 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5659 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5660 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5661 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5662 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5663 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5664 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5665 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5666 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5667 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5668 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5669 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5670 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5671 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5672 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5673 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5674 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5675 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5676 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5677 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5678 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5679 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5680 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5681 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5682 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5683 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5684 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5685 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5686 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5687 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5688 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5689 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5690 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5691 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5692 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5693 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5694 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5695 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5696 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5697 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5698 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5699 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5700 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5701 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5702 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5703 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5704 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5705 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5706 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5707 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5708 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5709 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5710 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5711 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5712 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5713 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5714 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5715 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5716 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5717 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5718 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5719 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5720 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5721 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5722 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5723 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5724 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5725 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5726 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5727 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5728 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5729 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5730 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5731 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5732 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5733 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5734 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5735 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5736 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5737 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5738 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5739 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5740 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5741 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5742 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5743 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5744 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5745 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5746 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5747 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5748 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5749 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5750 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5751 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5752 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5753 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5754 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5755 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5756 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5757 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5758 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5759 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5760 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5761 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5762 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5763 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5764 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5765 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5766 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5767 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5768 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5769 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5770 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5771 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5772 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5773 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5774 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5775 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5776 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5777 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5778 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5779 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5780 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5781 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5782 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5783 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5784 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5785 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5786 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5787 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5788 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5789 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5790 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5791 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5792 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5793 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5794 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5795 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5796 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5797 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5798 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5799 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5800 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5801 \$5373 \$5472 \$5372 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5802 \$5347 \$5472 \$5373 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5803 \$5374 \$5023 \$5347 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5804 \$5271 \$5023 \$5374 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5805 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5806 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5807 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5808 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5809 \$5376 \$5271 \$5375 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5810 \$5472 \$5271 \$5376 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5811 \$5377 \$5271 \$5472 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5812 \$5482 \$5271 \$5377 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5813 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5814 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5815 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5816 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5817 \$5378 \$5473 \$5473 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5818 AVDD|AVSS|VDD|VSS \$5473 \$5378 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5819 \$5379 \$5473 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5820 \$6150 \$5473 \$5379 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5821 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5822 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5823 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5824 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5825 \$5381 \$5474 \$5380 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5826 \$5348 \$5474 \$5381 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5827 \$5382 \$5027 \$5348 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5828 \$5272 \$5027 \$5382 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5829 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5830 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5831 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5832 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5833 \$5384 \$5272 \$5383 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5834 \$5474 \$5272 \$5384 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5835 \$5385 \$5272 \$5474 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5836 \$5483 \$5272 \$5385 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5837 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5838 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5839 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5840 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5841 \$5386 \$5475 \$5475 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5842 AVDD|AVSS|VDD|VSS \$5475 \$5386 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5843 \$5387 \$5475 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5844 \$6151 \$5475 \$5387 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5845 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5846 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5847 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5848 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5849 \$5389 \$5476 \$5388 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5850 \$5349 \$5476 \$5389 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5851 \$5390 \$5031 \$5349 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5852 \$5273 \$5031 \$5390 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5853 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5854 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5855 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5856 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5857 \$5392 \$5273 \$5391 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5858 \$5476 \$5273 \$5392 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5859 \$5393 \$5273 \$5476 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5860 \$5484 \$5273 \$5393 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5861 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5862 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5863 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5864 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5865 \$5394 \$5477 \$5477 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5866 AVDD|AVSS|VDD|VSS \$5477 \$5394 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5867 \$5395 \$5477 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5868 \$6152 \$5477 \$5395 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5869 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5870 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5871 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5872 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5873 \$5397 \$5478 \$5396 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5874 \$5350 \$5478 \$5397 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5875 \$5398 \$3346 \$5350 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5876 \$5274 \$3346 \$5398 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5877 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5878 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5879 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5880 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5881 \$5400 \$5274 \$5399 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5882 \$5478 \$5274 \$5400 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5883 \$5401 \$5274 \$5478 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5884 \$5485 \$5274 \$5401 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5885 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5886 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5887 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5888 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5889 \$5402 \$5479 \$5479 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5890 AVDD|AVSS|VDD|VSS \$5479 \$5402 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5891 \$5403 \$5479 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5892 \$6153 \$5479 \$5403 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5893 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5894 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5895 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5896 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5897 \$5405 \$5480 \$5404 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5898 \$5351 \$5480 \$5405 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5899 \$5406 \$3350 \$5351 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5900 \$5275 \$3350 \$5406 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5901 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5902 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5903 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5904 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5905 \$5408 \$5275 \$5407 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5906 \$5480 \$5275 \$5408 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5907 \$5409 \$5275 \$5480 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5908 \$5486 \$5275 \$5409 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5909 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5910 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5911 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5912 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5913 \$5410 \$5481 \$5481 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5914 AVDD|AVSS|VDD|VSS \$5481 \$5410 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5915 \$5411 \$5481 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5916 \$6154 \$5481 \$5411 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5917 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5918 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5919 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5920 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5921 \$5542 \$5023 \$5271 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5922 \$5347 \$5023 \$5542 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5923 \$5543 \$5472 \$5347 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5924 \$5372 \$5472 \$5543 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5925 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5926 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5927 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5928 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5929 \$5544 \$5271 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5930 \$5023 \$5271 \$5544 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5931 \$5545 \$5271 \$5023 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5932 AVDD|AVSS|VDD|VSS \$5271 \$5545 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5933 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5934 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5935 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5936 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5937 \$5546 \$5473 \$6150 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5938 AVDD|AVSS|VDD|VSS \$5473 \$5546 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5939 \$5547 \$5473 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5940 \$5473 \$5473 \$5547 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5941 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5942 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5943 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5944 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5945 \$5548 \$5027 \$5272 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5946 \$5348 \$5027 \$5548 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5947 \$5549 \$5474 \$5348 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5948 \$5380 \$5474 \$5549 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5949 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5950 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5951 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5952 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5953 \$5550 \$5272 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5954 \$5027 \$5272 \$5550 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5955 \$5551 \$5272 \$5027 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5956 AVDD|AVSS|VDD|VSS \$5272 \$5551 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5957 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5958 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5959 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5960 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5961 \$5552 \$5475 \$6151 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5962 AVDD|AVSS|VDD|VSS \$5475 \$5552 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5963 \$5553 \$5475 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5964 \$5475 \$5475 \$5553 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5965 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5966 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5967 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5968 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5969 \$5554 \$5031 \$5273 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5970 \$5349 \$5031 \$5554 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5971 \$5555 \$5476 \$5349 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5972 \$5388 \$5476 \$5555 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5973 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5974 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5975 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5976 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5977 \$5556 \$5273 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5978 \$5031 \$5273 \$5556 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5979 \$5557 \$5273 \$5031 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5980 AVDD|AVSS|VDD|VSS \$5273 \$5557 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5981 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5982 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5983 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5984 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5985 \$5558 \$5477 \$6152 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5986 AVDD|AVSS|VDD|VSS \$5477 \$5558 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$5987 \$5559 \$5477 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5988 \$5477 \$5477 \$5559 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5989 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5990 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5991 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5992 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5993 \$5560 \$3346 \$5274 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5994 \$5350 \$3346 \$5560 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5995 \$5561 \$5478 \$5350 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$5996 \$5396 \$5478 \$5561 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$5997 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5998 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5999 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6000 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6001 \$5562 \$5274 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6002 \$3346 \$5274 \$5562 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6003 \$5563 \$5274 \$3346 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6004 AVDD|AVSS|VDD|VSS \$5274 \$5563 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6005 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6006 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6007 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6008 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6009 \$5564 \$5479 \$6153 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6010 AVDD|AVSS|VDD|VSS \$5479 \$5564 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6011 \$5565 \$5479 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6012 \$5479 \$5479 \$5565 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6013 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6014 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6015 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6016 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6017 \$5566 \$3350 \$5275 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6018 \$5351 \$3350 \$5566 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6019 \$5567 \$5480 \$5351 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6020 \$5404 \$5480 \$5567 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6021 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6022 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6023 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6024 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6025 \$5568 \$5275 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6026 \$3350 \$5275 \$5568 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6027 \$5569 \$5275 \$3350 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6028 AVDD|AVSS|VDD|VSS \$5275 \$5569 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6029 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6030 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6031 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6032 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6033 \$5570 \$5481 \$6154 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6034 AVDD|AVSS|VDD|VSS \$5481 \$5570 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6035 \$5571 \$5481 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6036 \$5481 \$5481 \$5571 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6037 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6038 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6039 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6040 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6041 \$5677 \$5472 \$5372 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6042 \$5347 \$5472 \$5677 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6043 \$5678 \$5023 \$5347 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6044 \$5271 \$5023 \$5678 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6045 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6046 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6047 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6048 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6049 \$5679 \$5271 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6050 \$5023 \$5271 \$5679 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6051 \$5680 \$5271 \$5023 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6052 AVDD|AVSS|VDD|VSS \$5271 \$5680 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6053 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6054 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6055 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6056 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6057 \$5681 \$5473 \$5473 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6058 AVDD|AVSS|VDD|VSS \$5473 \$5681 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6059 \$5682 \$5473 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6060 \$6150 \$5473 \$5682 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6061 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6062 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6063 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6064 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6065 \$5683 \$5474 \$5380 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6066 \$5348 \$5474 \$5683 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6067 \$5684 \$5027 \$5348 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6068 \$5272 \$5027 \$5684 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6069 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6070 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6071 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6072 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6073 \$5685 \$5272 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6074 \$5027 \$5272 \$5685 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6075 \$5686 \$5272 \$5027 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6076 AVDD|AVSS|VDD|VSS \$5272 \$5686 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6077 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6078 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6079 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6080 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6081 \$5687 \$5475 \$5475 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6082 AVDD|AVSS|VDD|VSS \$5475 \$5687 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6083 \$5688 \$5475 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6084 \$6151 \$5475 \$5688 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6085 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6086 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6087 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6088 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6089 \$5689 \$5476 \$5388 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6090 \$5349 \$5476 \$5689 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6091 \$5690 \$5031 \$5349 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6092 \$5273 \$5031 \$5690 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6093 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6094 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6095 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6096 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6097 \$5691 \$5273 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6098 \$5031 \$5273 \$5691 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6099 \$5692 \$5273 \$5031 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6100 AVDD|AVSS|VDD|VSS \$5273 \$5692 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6101 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6102 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6103 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6104 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6105 \$5693 \$5477 \$5477 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6106 AVDD|AVSS|VDD|VSS \$5477 \$5693 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6107 \$5694 \$5477 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6108 \$6152 \$5477 \$5694 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6109 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6110 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6111 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6112 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6113 \$5695 \$5478 \$5396 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6114 \$5350 \$5478 \$5695 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6115 \$5696 \$3346 \$5350 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6116 \$5274 \$3346 \$5696 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6117 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6118 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6119 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6120 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6121 \$5697 \$5274 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6122 \$3346 \$5274 \$5697 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6123 \$5698 \$5274 \$3346 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6124 AVDD|AVSS|VDD|VSS \$5274 \$5698 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6125 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6126 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6127 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6128 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6129 \$5699 \$5479 \$5479 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6130 AVDD|AVSS|VDD|VSS \$5479 \$5699 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6131 \$5700 \$5479 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6132 \$6153 \$5479 \$5700 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6133 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6134 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6135 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6136 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6137 \$5701 \$5480 \$5404 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6138 \$5351 \$5480 \$5701 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6139 \$5702 \$3350 \$5351 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6140 \$5275 \$3350 \$5702 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6141 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6142 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6143 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6144 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6145 \$5703 \$5275 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6146 \$3350 \$5275 \$5703 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6147 \$5704 \$5275 \$3350 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6148 AVDD|AVSS|VDD|VSS \$5275 \$5704 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6149 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6150 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6151 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6152 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6153 \$5705 \$5481 \$5481 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6154 AVDD|AVSS|VDD|VSS \$5481 \$5705 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6155 \$5706 \$5481 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6156 \$6154 \$5481 \$5706 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6157 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6158 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6159 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6160 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6161 \$5822 \$5023 \$5271 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6162 \$5347 \$5023 \$5822 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6163 \$5823 \$5472 \$5347 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6164 \$5372 \$5472 \$5823 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6165 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6166 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6167 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6168 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6169 \$5824 \$5271 \$5482 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6170 \$5472 \$5271 \$5824 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6171 \$5825 \$5271 \$5472 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6172 \$5375 \$5271 \$5825 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6173 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6174 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6175 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6176 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6177 \$5826 \$5473 \$6150 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6178 AVDD|AVSS|VDD|VSS \$5473 \$5826 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6179 \$5827 \$5473 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6180 \$5473 \$5473 \$5827 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6181 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6182 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6183 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6184 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6185 \$5828 \$5027 \$5272 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6186 \$5348 \$5027 \$5828 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6187 \$5829 \$5474 \$5348 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6188 \$5380 \$5474 \$5829 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6189 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6190 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6191 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6192 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6193 \$5830 \$5272 \$5483 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6194 \$5474 \$5272 \$5830 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6195 \$5831 \$5272 \$5474 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6196 \$5383 \$5272 \$5831 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6197 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6198 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6199 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6200 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6201 \$5832 \$5475 \$6151 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6202 AVDD|AVSS|VDD|VSS \$5475 \$5832 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6203 \$5833 \$5475 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6204 \$5475 \$5475 \$5833 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6205 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6206 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6207 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6208 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6209 \$5834 \$5031 \$5273 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6210 \$5349 \$5031 \$5834 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6211 \$5835 \$5476 \$5349 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6212 \$5388 \$5476 \$5835 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6213 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6214 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6215 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6216 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6217 \$5836 \$5273 \$5484 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6218 \$5476 \$5273 \$5836 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6219 \$5837 \$5273 \$5476 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6220 \$5391 \$5273 \$5837 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6221 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6222 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6223 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6224 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6225 \$5838 \$5477 \$6152 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6226 AVDD|AVSS|VDD|VSS \$5477 \$5838 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6227 \$5839 \$5477 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6228 \$5477 \$5477 \$5839 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6229 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6230 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6231 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6232 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6233 \$5840 \$3346 \$5274 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6234 \$5350 \$3346 \$5840 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6235 \$5841 \$5478 \$5350 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6236 \$5396 \$5478 \$5841 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6237 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6238 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6239 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6240 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6241 \$5842 \$5274 \$5485 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6242 \$5478 \$5274 \$5842 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6243 \$5843 \$5274 \$5478 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6244 \$5399 \$5274 \$5843 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6245 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6246 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6247 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6248 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6249 \$5844 \$5479 \$6153 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6250 AVDD|AVSS|VDD|VSS \$5479 \$5844 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6251 \$5845 \$5479 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6252 \$5479 \$5479 \$5845 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6253 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6254 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6255 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6256 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6257 \$5846 \$3350 \$5275 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6258 \$5351 \$3350 \$5846 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6259 \$5847 \$5480 \$5351 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6260 \$5404 \$5480 \$5847 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6261 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6262 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6263 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6264 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6265 \$5848 \$5275 \$5486 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6266 \$5480 \$5275 \$5848 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6267 \$5849 \$5275 \$5480 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6268 \$5407 \$5275 \$5849 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6269 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6270 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6271 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6272 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6273 \$5850 \$5481 \$6154 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6274 AVDD|AVSS|VDD|VSS \$5481 \$5850 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6275 \$5851 \$5481 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6276 \$5481 \$5481 \$5851 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6277 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6278 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6279 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6280 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6281 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6282 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6283 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6284 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6285 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6286 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6287 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6288 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6289 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6290 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6291 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6292 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6293 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6294 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6295 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6296 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6297 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6298 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6299 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6300 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6301 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6302 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6303 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6304 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6305 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6306 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6307 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6308 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6309 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6310 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6311 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6312 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6313 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6314 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6315 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6316 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6317 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6318 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6319 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6320 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6321 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6322 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6323 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6324 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6325 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6326 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6327 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6328 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6329 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6330 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6331 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6332 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6333 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6334 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6335 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6336 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6337 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6338 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6339 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6340 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6341 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6342 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6343 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6344 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6345 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6346 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6347 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6348 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6349 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6350 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6351 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6352 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6353 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6354 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6355 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6356 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6357 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6358 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6359 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6360 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6361 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6362 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6363 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6364 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6365 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6366 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6367 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6368 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6369 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6370 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6371 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6372 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6373 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6374 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6375 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6376 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6377 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6378 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6379 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6380 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6381 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6382 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6383 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6384 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6385 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6386 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6387 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6388 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6389 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6390 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6391 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6392 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6393 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6394 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6395 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6396 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6397 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6398 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6399 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6400 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6401 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6402 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6403 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6404 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6405 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6406 ISBCS2 ISBCS2 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=6U W=2U
+ AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6407 \$6841 ISBCS2 \$6811 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$6408 \$6795 ISBCS2 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=6U W=2U
+ AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6409 \$6795 ISBCS2 \$6811 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$6410 \$6841 ISBCS2 \$7527 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$6411 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6412 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6413 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6414 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6415 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6416 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6417 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U PD=5.72U
M$6418 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U PD=5.72U
M$6419 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U PD=5.72U
M$6420 AVDD|AVSS|VDD|VSS \$6812 \$6797 gf180mcu_gnd nfet_03v3 L=2U W=2.25U
+ AS=1.3725P AD=0.9P PS=5.72U PD=3.05U
M$6421 \$6797 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2.25U
+ AS=0.9P AD=1.3725P PS=3.05U PD=5.72U
M$6422 AVDD|AVSS|VDD|VSS \$6812 \$6812 gf180mcu_gnd nfet_03v3 L=2U W=2.25U
+ AS=1.3725P AD=0.9P PS=5.72U PD=3.05U
M$6423 \$6812 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2.25U
+ AS=0.9P AD=1.3725P PS=3.05U PD=5.72U
M$6424 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U PD=3.05U
M$6425 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U PD=5.72U
M$6426 AVDD|AVSS|VDD|VSS \$6812 \$6812 gf180mcu_gnd nfet_03v3 L=2U W=2.25U
+ AS=1.3725P AD=0.9P PS=5.72U PD=3.05U
M$6427 \$6812 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2.25U
+ AS=0.9P AD=1.3725P PS=3.05U PD=5.72U
M$6428 AVDD|AVSS|VDD|VSS \$6812 \$6797 gf180mcu_gnd nfet_03v3 L=2U W=2.25U
+ AS=1.3725P AD=0.9P PS=5.72U PD=3.05U
M$6429 \$6797 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2.25U
+ AS=0.9P AD=1.3725P PS=3.05U PD=5.72U
M$6430 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U PD=3.05U
M$6431 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U PD=5.72U
M$6432 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U PD=5.72U
M$6433 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U PD=5.72U
M$6434 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U PD=5.72U
M$6435 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U PD=3.62U
M$6436 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U PD=3.62U
M$6437 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U PD=3.62U
M$6438 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U PD=3.62U
M$6439 \$6844 \$6843 \$6842 gf180mcu_gnd nfet_03v3 L=2U W=1.2U AS=0.732P
+ AD=0.48P PS=3.62U PD=2U
M$6440 AVDD|AVSS|VDD|VSS \$6843 \$6844 gf180mcu_gnd nfet_03v3 L=2U W=1.2U
+ AS=0.48P AD=0.732P PS=2U PD=3.62U
M$6441 \$7258 \$6843 \$6842 gf180mcu_gnd nfet_03v3 L=2U W=1.2U AS=0.732P
+ AD=0.48P PS=3.62U PD=2U
M$6442 \$7259 \$6843 \$7258 gf180mcu_gnd nfet_03v3 L=2U W=1.2U AS=0.48P
+ AD=0.732P PS=2U PD=3.62U
M$6443 \$7800 \$6843 \$6843 gf180mcu_gnd nfet_03v3 L=2U W=1.2U AS=0.732P
+ AD=0.48P PS=3.62U PD=2U
M$6444 \$7259 \$6843 \$7800 gf180mcu_gnd nfet_03v3 L=2U W=1.2U AS=0.48P
+ AD=0.732P PS=2U PD=3.62U
M$6445 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P PS=3.62U PD=2U
M$6446 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U PD=3.62U
M$6447 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U PD=3.62U
M$6448 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U PD=3.62U
M$6449 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U PD=3.62U
M$6450 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U PD=3.62U
M$6451 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6452 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6453 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6454 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6455 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6456 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6457 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6458 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6459 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6460 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6461 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6462 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6463 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6464 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6465 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6466 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6467 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6468 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6469 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6470 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6471 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6472 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6473 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6474 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6475 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6476 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6477 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6478 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6479 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6480 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6481 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6482 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6483 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6484 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6485 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6486 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6487 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6488 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6489 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6490 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6491 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6492 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6493 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6494 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6495 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6496 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6497 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6498 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6499 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6500 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6501 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6502 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6503 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6504 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6505 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6506 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6507 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6508 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6509 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6510 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6511 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6512 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6513 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6514 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6515 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6516 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6517 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6518 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6519 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6520 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6521 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6522 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6523 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6524 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6525 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6526 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6527 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6528 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6529 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6530 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6531 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6532 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6533 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6534 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6535 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6536 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6537 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6538 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6539 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6540 IREF ISBCS2 \$7527 gf180mcu_gnd nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$6541 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6542 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U PD=5.72U
M$6543 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U PD=3.05U
M$6544 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U PD=5.72U
M$6545 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U PD=3.05U
M$6546 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U PD=5.72U
M$6547 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U PD=5.72U
M$6548 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U PD=3.62U
M$6549 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P PS=3.62U PD=2U
M$6550 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U PD=3.62U
M$6551 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U PD=3.62U
M$6552 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6553 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6554 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6555 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6556 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6557 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6558 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6559 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6560 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6561 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6562 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6563 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6564 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6565 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6566 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6567 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6568 AVDD|AVSS|VDD|VSS \$6812 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6569 \$6762 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6570 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U
+ AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6571 \$6793 \$6812 AVDD|AVSS|VDD|VSS gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=0.8P PS=2.8U PD=2.8U
M$6572 AVDD|AVSS|VDD|VSS \$6812 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P
+ AD=1.22P PS=2.8U PD=5.22U
M$6573 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6574 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6575 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6576 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6577 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6578 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6579 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6580 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6581 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6582 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6583 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6584 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6585 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6586 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6587 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6588 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6589 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6590 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6591 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6592 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6593 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6594 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6595 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6596 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6597 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6598 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6599 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6600 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6601 \$12262 \$6843 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6602 \$6793 \$6843 \$12262 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P
+ PS=2.8U PD=2.8U
M$6603 \$12262 \$6843 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6604 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6605 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6606 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6607 \$6762 \$6843 B1|VOUT gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6608 B1|VOUT \$6843 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P
+ PS=2.8U PD=2.8U
M$6609 \$6762 \$6843 B1|VOUT gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6610 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6611 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6612 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6613 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6614 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6615 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6616 \$12262 \$6843 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6617 \$6793 \$6843 \$12262 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P
+ PS=2.8U PD=2.8U
M$6618 \$12262 \$6843 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6619 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6620 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6621 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6622 B1|VOUT \$6843 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6623 \$6762 \$6843 B1|VOUT gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P
+ PS=2.8U PD=2.8U
M$6624 B1|VOUT \$6843 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6625 \$12262 \$6843 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6626 \$6793 \$6843 \$12262 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P
+ PS=2.8U PD=2.8U
M$6627 \$12262 \$6843 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6628 \$6762 \$6843 B1|VOUT gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6629 B1|VOUT \$6843 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P
+ PS=2.8U PD=2.8U
M$6630 \$6762 \$6843 B1|VOUT gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6631 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6632 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6633 B1|VOUT \$6843 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6634 \$6762 \$6843 B1|VOUT gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P
+ PS=2.8U PD=2.8U
M$6635 B1|VOUT \$6843 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6636 \$12262 \$6843 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6637 \$6793 \$6843 \$12262 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P
+ PS=2.8U PD=2.8U
M$6638 \$12262 \$6843 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6639 \$6762 \$6843 B1|VOUT gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6640 B1|VOUT \$6843 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P
+ PS=2.8U PD=2.8U
M$6641 \$6762 \$6843 B1|VOUT gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6642 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6643 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6644 \$12262 \$6843 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6645 \$6793 \$6843 \$12262 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P
+ PS=2.8U PD=2.8U
M$6646 \$12262 \$6843 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6647 B1|VOUT \$6843 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6648 \$6762 \$6843 B1|VOUT gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P
+ PS=2.8U PD=2.8U
M$6649 B1|VOUT \$6843 \$6762 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6650 \$6793 \$6843 \$12262 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P
+ PS=5.22U PD=2.8U
M$6651 \$12262 \$6843 \$6793 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P
+ PS=2.8U PD=2.8U
M$6652 \$6793 \$6843 \$12262 gf180mcu_gnd nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P
+ PS=2.8U PD=5.22U
M$6653 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6654 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6655 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6656 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6657 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6658 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6659 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6660 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6661 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6662 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6663 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6664 AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS AVDD|AVSS|VDD|VSS gf180mcu_gnd
+ nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
C$6665 \$2476 \$2575 1.9208e-13 cap_mim_2f0_m4m5_noshield A=96.04P P=39.2U
C$6666 A1|VN B1|VOUT 1.9208e-13 cap_mim_2f0_m4m5_noshield A=96.04P P=39.2U
C$6667 \$6832 \$6833 2e-11 cap_mim_2f0_m4m5_noshield A=10000P P=400U
C$6668 \$24461 \$24462 2e-11 cap_mim_2f0_m4m5_noshield A=10000P P=400U
.ENDS Filter_TOP
