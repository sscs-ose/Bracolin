* Extracted by KLayout with GF180MCU LVS runset on : 25/04/2024 15:23

.SUBCKT track_Dyn VSSA clks Vinp Vinn Vcom VDP VDN CK1 vocp VDDD A B C
M$1 \$13 clks \$45 \$45 pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$2 \$14 \$13 \$45 \$45 pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$3 \$45 \$49 \$183 \$183 pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U PD=9.3U
M$4 \$49 \$17 \$183 \$183 pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U PD=9.3U
M$5 \$185 \$22 \$20 \$185 pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U PD=9.3U
M$6 \$185 \$20 \$45 \$185 pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U PD=9.3U
M$7 \$1126 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$8 \$1127 CK1 \$1126 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$9 \$1064 \$1063 \$1127 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$10 \$1076 \$1064 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$11 \$17 \$14 \$45 \$45 pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U PD=9.3U
M$12 \$45 \$14 \$22 \$45 pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U PD=9.3U
M$13 \$1070 \$1076 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$14 \$1107 \$1070 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$15 \$1109 \$1108 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$16 vocp \$1083 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$17 \$1168 \$1179 \$1108 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$18 \$1108 \$1179 \$1168 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$19 \$1168 \$1179 \$1108 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$20 \$1108 \$1179 \$1168 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$21 \$1169 \$1101 \$1083 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$22 \$1083 \$1101 \$1169 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$23 \$1169 \$1101 \$1083 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$24 \$1083 \$1101 \$1169 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$25 \$1179 \$1070 VDDD VDDD pfet_03v3 L=0.28U W=2.35U AS=1.5275P AD=1.5275P
+ PS=6U PD=6U
M$26 VDDD \$1070 \$1179 VDDD pfet_03v3 L=0.28U W=2.35U AS=1.5275P AD=1.5275P
+ PS=6U PD=6U
M$27 \$1101 \$1070 VDDD VDDD pfet_03v3 L=0.28U W=2.35U AS=1.5275P AD=1.5275P
+ PS=6U PD=6U
M$28 VDDD \$1070 \$1101 VDDD pfet_03v3 L=0.28U W=2.35U AS=1.5275P AD=1.5275P
+ PS=6U PD=6U
M$29 VDDD \$1083 \$1168 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$30 \$1168 \$1083 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$31 VDDD \$1083 \$1168 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$32 \$1168 \$1083 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$33 VDDD \$1108 \$1169 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$34 \$1169 \$1108 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$35 VDDD \$1108 \$1169 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$36 \$1169 \$1108 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$37 \$1063 vocp VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$38 VDDD \$1109 \$1063 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$39 \$13 clks VSSA VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$40 \$14 \$13 VSSA VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$41 VDP VSSA Vcom VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$42 VDP \$49 Vinp VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$43 VDP VSSA Vcom VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$44 VDP \$49 Vinp VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$45 VDP VSSA Vcom VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$46 VDP \$49 Vinp VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$47 VDP VSSA Vcom VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$48 VDP \$49 Vinp VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$49 VDP VSSA Vcom VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$50 VDP \$49 Vinp VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$51 \$17 \$14 \$16 VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$52 \$17 \$49 \$16 VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$53 VSSA \$13 \$16 VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$54 Vinp \$49 \$16 VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$55 \$18 \$45 \$49 VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$56 VSSA \$13 \$18 VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$57 \$19 \$13 VSSA VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$58 \$20 \$45 \$19 VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$59 \$21 \$20 Vinn VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$60 \$21 \$13 VSSA VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$61 \$21 \$20 \$22 VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$62 \$21 \$14 \$22 VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$63 Vinn \$20 VDN VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$64 Vcom VSSA VDN VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$65 Vinn \$20 VDN VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$66 Vcom VSSA VDN VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$67 Vinn \$20 VDN VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$68 Vcom VSSA VDN VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$69 Vinn \$20 VDN VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$70 Vcom VSSA VDN VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$71 Vinn \$20 VDN VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$72 Vcom VSSA VDN VSSA nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$73 \$1064 clks VSSA VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$74 VSSA CK1 \$1064 VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$75 VSSA \$1063 \$1064 VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$76 \$1068 \$1064 \$1076 VSSA nfet_03v3 L=35U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$77 \$1068 \$1064 VSSA VSSA nfet_03v3 L=35U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$78 \$1098 \$1064 \$1128 VSSA nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$79 \$1076 A \$1128 VSSA nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$80 \$1098 \$1064 VSSA VSSA nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$81 \$1099 \$1064 \$1129 VSSA nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$82 \$1099 \$1064 VSSA VSSA nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$83 \$1076 B \$1129 VSSA nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$84 \$1100 \$1064 VSSA VSSA nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$85 \$1100 \$1064 \$1130 VSSA nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$86 \$1076 C \$1130 VSSA nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$87 \$1070 \$1076 VSSA VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$88 \$1114 VDP \$1101 VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$89 \$1114 VDN \$1179 VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$90 \$1179 VDN \$1114 VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$91 \$1101 VDP \$1114 VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$92 \$1114 \$1070 VSSA VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$93 \$1114 VDP \$1101 VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$94 \$1114 VDN \$1179 VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$95 VSSA \$1070 \$1114 VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$96 \$1179 VDN \$1114 VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$97 \$1101 VDP \$1114 VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$98 \$1114 \$1070 VSSA VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$99 \$1114 VDP \$1101 VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$100 \$1114 VDN \$1179 VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$101 \$1101 VDP \$1114 VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$102 \$1179 VDN \$1114 VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$103 \$1107 \$1070 VSSA VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$104 \$1108 \$1107 VSSA VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$105 VSSA \$1108 \$1083 VSSA nfet_03v3 L=0.28U W=6.3U AS=3.843P AD=2.52P
+ PS=13.82U PD=7.1U
M$106 \$1108 \$1083 VSSA VSSA nfet_03v3 L=0.28U W=6.3U AS=2.52P AD=3.843P
+ PS=7.1U PD=13.82U
M$107 \$1083 \$1107 VSSA VSSA nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$108 \$1109 \$1108 VSSA VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$109 vocp \$1083 VSSA VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$110 \$1085 vocp VSSA VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$111 \$1063 \$1109 \$1085 VSSA nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
C$112 \$16 \$183 2e-13 cap_mim_2f0_m4m5_noshield A=100P P=40U
C$113 \$16 \$183 2e-13 cap_mim_2f0_m4m5_noshield A=100P P=40U
C$114 \$16 \$183 2e-13 cap_mim_2f0_m4m5_noshield A=100P P=40U
C$115 \$21 \$185 2e-13 cap_mim_2f0_m4m5_noshield A=100P P=40U
C$116 \$21 \$185 2e-13 cap_mim_2f0_m4m5_noshield A=100P P=40U
C$117 \$21 \$185 2e-13 cap_mim_2f0_m4m5_noshield A=100P P=40U
.ENDS track_Dyn
