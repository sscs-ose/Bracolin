* Extracted by KLayout with GF180MCU LVS runset on : 04/01/2024 18:11

.SUBCKT CM_iref ISBCS2 IREF VSS
M$1 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$2 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$3 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5 ISBCS2 ISBCS2 VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$7 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$8 \$13 ISBCS2 VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$9 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$10 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$11 \$13 ISBCS2 \$19 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$12 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$13 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$14 \$24 ISBCS2 \$19 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$15 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$16 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$17 \$24 ISBCS2 \$31 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$18 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$19 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$20 IREF ISBCS2 \$31 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$21 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$22 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$23 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$24 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
.ENDS CM_iref
