* NGSPICE file created from PRbiased_net.ext - technology: gf180mcuD

.subckt PRbiased_net VSS VDD ITN IBN VA IBP VB ITP
X0 ITP IBP.t4 a_12130_9713# VDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1 a_412_1806# IBN.t4 a_n160_7781.t3 VSS.t19 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2 VSS.t225 VSS.t224 VSS.t225 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3 VDD.t222 VDD.t221 VDD.t222 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4 VDD.t220 VDD.t219 VDD.t220 VDD.t80 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5 VSS.t223 VSS.t222 VSS.t223 VSS.t29 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6 a_12101_2572# a_11579_648.t5 a_11579_648.t6 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X7 a_6218_1806# a_n160_7781.t8 VDD.t226 VSS.t6 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X8 VDD.t218 VDD.t217 VDD.t218 VDD.t24 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X9 VDD.t216 VDD.t215 VDD.t216 VDD.t24 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X10 a_1776_9713# a_n160_6615.t13 VDD.t224 VDD.t15 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X11 VDD.t214 VDD.t213 VDD.t214 VDD.t142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X12 VSS.t221 VSS.t220 VSS.t221 VSS.t18 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X13 VSS.t219 VSS.t218 VSS.t219 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X14 VDD.t212 VDD.t211 VDD.t212 VDD.t21 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X15 ITP a_12_588.t3 a_12130_8547# VDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X16 VSS.t217 VSS.t216 VSS.t217 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X17 VSS.t215 VSS.t214 VSS.t215 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X18 VSS.t213 VSS.t212 VSS.t213 VSS.t3 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X19 VDD.t210 VDD.t209 VDD.t210 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X20 ITP a_12_588.t3 a_12130_6615# VDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X21 VSS.t211 VSS.t210 VSS.t211 VSS.t49 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X22 VDD.t208 VDD.t207 VDD.t208 VDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X23 VDD.t206 VDD.t205 VDD.t206 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X24 VDD.t204 VDD.t203 VDD.t204 VDD.t80 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X25 VDD.t202 VDD.t201 VDD.t202 VDD.t80 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X26 VSS.t209 VSS.t208 VSS.t209 VSS.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X27 VSS.t207 VSS.t206 VSS.t207 VSS.t32 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X28 VDD.t200 VDD.t199 VDD.t200 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X29 VDD.t198 VDD.t197 VDD.t198 VDD.t24 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X30 VSS.t205 VSS.t204 VSS.t205 VSS.t59 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X31 a_1776_8547# a_n160_6615.t16 VDD.t16 VDD.t15 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X32 VDD.t196 VDD.t195 VDD.t196 VDD.t142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X33 a_1776_6615# a_n160_6615.t17 VDD.t17 VDD.t15 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X34 VDD.t194 VDD.t193 VDD.t194 VDD.t142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X35 a_1816_3730# a_12_588.t2 ITN.t5 VSS.t20 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X36 VSS.t203 VSS.t202 VSS.t203 VSS.t41 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X37 VSS.t201 VSS.t200 VSS.t201 VSS.t38 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X38 a_13505_3730# a_11579_648.t12 VSS.t9 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X39 VDD.t192 VDD.t191 VDD.t192 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X40 VSS.t199 VSS.t198 VSS.t199 VSS.t1 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X41 VDD.t190 VDD.t189 VDD.t190 VDD.t2 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X42 VDD.t188 VDD.t187 VDD.t188 VDD.t8 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X43 VSS.t197 VSS.t196 VSS.t197 VSS.t46 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X44 VDD.t186 VDD.t185 VDD.t186 VDD.t149 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X45 VDD.t184 VDD.t183 VDD.t184 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X46 VDD.t182 VDD.t181 VDD.t182 VDD.t80 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X47 VSS.t195 VSS.t194 VSS.t195 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X48 VDD.t180 VDD.t179 VDD.t180 VDD.t24 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X49 VDD.t178 VDD.t177 VDD.t178 VDD.t75 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X50 VDD.t176 VDD.t175 VDD.t176 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X51 VDD.t174 VDD.t173 VDD.t174 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X52 a_1816_648# IBN.t6 ITN.t2 VSS.t20 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X53 a_12101_648# a_11579_648.t9 a_11579_648.t10 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X54 VDD.t172 VDD.t171 VDD.t172 VDD.t15 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X55 VDD.t170 VDD.t169 VDD.t170 VDD.t100 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X56 VDD.t168 VDD.t167 VDD.t168 VDD.t142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X57 VSS.t193 VSS.t192 VSS.t193 VSS.t59 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X58 VSS.t191 VSS.t190 VSS.t191 VSS.t26 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X59 VSS.t189 VSS.t188 VSS.t189 VSS.t23 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X60 ITP IBP.t5 a_12130_7781# VDD.t8 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X61 VSS a_11579_648.t14 a_12101_3730# VSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X62 VDD.t166 VDD.t165 VDD.t166 VDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X63 VDD.t164 VDD.t163 VDD.t164 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X64 a_13505_648# a_11579_648.t15 VSS.t230 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X65 VDD.t162 VDD.t161 VDD.t162 VDD.t37 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X66 VDD.t160 VDD.t159 VDD.t160 VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X67 VDD.t158 VDD.t157 VDD.t158 VDD.t80 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X68 VDD.t156 VDD.t155 VDD.t156 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X69 a_1816_2572# IBN.t8 ITN.t0 VSS.t20 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X70 a_13505_2572# a_11579_648.t17 VSS.t8 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X71 a_412_3730# IBN.t9 a_n160_7781.t1 VSS.t19 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X72 VSS.t187 VSS.t186 VSS.t187 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X73 VSS.t185 VSS.t184 VSS.t185 VSS.t46 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X74 VSS.t183 VSS.t182 VSS.t183 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X75 VSS.t181 VSS.t180 VSS.t181 VSS.t3 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X76 VSS.t179 VSS.t178 VSS.t179 VSS.t29 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X77 a_1776_7781# a_n160_6615.t19 VDD.t227 VDD.t15 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X78 VDD.t154 VDD.t153 VDD.t154 VDD.t142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X79 VDD.t152 VDD.t151 VDD.t152 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X80 VDD.t150 VDD.t148 VDD.t150 VDD.t149 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X81 VA a_5850_6555.t8 a_7656_9713# VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X82 VDD.t147 VDD.t146 VDD.t147 VDD.t75 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X83 VSS.t177 VSS.t176 VSS.t177 VSS.t32 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X84 a_6218_3730# a_n160_7781.t10 a_5696_3730.t0 VSS.t6 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X85 ITN IBN.t10 a_412_1806# VSS.t18 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X86 VDD.t145 VDD.t144 VDD.t145 VDD.t100 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X87 VDD.t143 VDD.t141 VDD.t143 VDD.t142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X88 VDD.t140 VDD.t139 VDD.t140 VDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X89 VDD.t138 VDD.t137 VDD.t138 VDD.t100 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X90 VSS.t175 VSS.t174 VSS.t175 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X91 VDD.t136 VDD.t135 VDD.t136 VDD.t37 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X92 VDD.t134 VDD.t133 VDD.t134 VDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X93 VDD.t132 VDD.t131 VDD.t132 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X94 VSS.t173 VSS.t172 VSS.t173 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X95 VSS a_11579_648.t18 a_12101_2572# VSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X96 VDD.t130 VDD.t129 VDD.t130 VDD.t37 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X97 a_7656_9713# a_5850_6555.t9 a_5696_648.t2 VDD.t4 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X98 VDD.t128 VDD.t127 VDD.t128 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X99 VSS.t171 VSS.t170 VSS.t171 VSS.t49 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X100 VDD.t126 VDD.t125 VDD.t126 VDD.t100 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X101 VDD.t124 VDD.t122 VDD.t124 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X102 VSS.t169 VSS.t168 VSS.t169 VSS.t26 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X103 IBN a_n160_7781.t12 a_6218_1806# VSS.t5 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X104 VSS.t167 VSS.t166 VSS.t167 VSS.t1 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X105 VDD.t121 VDD.t120 VDD.t121 VDD.t7 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X106 a_412_2572# a_12_588.t2 a_n160_6615.t10 VSS.t19 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X107 VSS.t165 VSS.t164 VSS.t165 VSS.t41 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X108 a_7622_648# a_n160_7781.t13 a_12_588.t2 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X109 VSS.t163 VSS.t162 VSS.t163 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X110 IBP a_5850_6555.t10 a_7656_8547# VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X111 VDD.t119 VDD.t118 VDD.t119 VDD.t75 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X112 VSS.t161 VSS.t160 VSS.t161 VSS.t59 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X113 VSS.t159 VSS.t158 VSS.t159 VSS.t23 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X114 VSS.t157 VSS.t156 VSS.t157 VSS.t29 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X115 VB a_5850_6555.t11 a_7656_6615# VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X116 VDD.t117 VDD.t116 VDD.t117 VDD.t75 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X117 VDD.t115 VDD.t114 VDD.t115 VDD.t40 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X118 VSS.t155 VSS.t154 VSS.t155 VSS.t21 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X119 a_6218_648# a_n160_7781.t14 a_5696_648.t0 VSS.t6 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X120 VDD.t113 VDD.t112 VDD.t113 VDD.t100 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X121 VSS.t153 VSS.t152 VSS.t153 VSS.t38 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X122 VSS.t151 VSS.t150 VSS.t151 VSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X123 a_6218_2572# a_n160_7781.t15 VDD.t225 VSS.t6 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X124 VSS.t149 VSS.t148 VSS.t149 VSS.t20 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X125 VSS.t147 VSS.t146 VSS.t147 VSS.t7 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X126 VDD.t111 VDD.t110 VDD.t111 VDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X127 VDD.t109 VDD.t108 VDD.t109 VDD.t37 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X128 a_7656_8547# a_5850_6555.t12 VSS.t10 VDD.t4 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X129 VDD.t107 VDD.t106 VDD.t107 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X130 VSS.t145 VSS.t144 VSS.t145 VSS.t41 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X131 VSS.t143 VSS.t142 VSS.t143 VSS.t38 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X132 VSS.t141 VSS.t140 VSS.t141 VSS.t46 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X133 a_7656_6615# a_5850_6555.t13 a_5696_3730.t2 VDD.t4 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X134 a_13536_9713# a_12_588.t3 ITP.t7 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X135 VDD.t105 VDD.t104 VDD.t105 VDD.t8 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X136 VDD.t103 VDD.t102 VDD.t103 VDD.t9 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X137 VDD.t101 VDD.t99 VDD.t101 VDD.t100 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X138 VDD.t98 VDD.t97 VDD.t98 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X139 VDD.t96 VDD.t95 VDD.t96 VDD.t75 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X140 VDD.t94 VDD.t92 VDD.t94 VDD.t93 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X141 VDD.t91 VDD.t90 VDD.t91 VDD.t37 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X142 VDD.t89 VDD.t88 VDD.t89 VDD.t40 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X143 VDD.t87 VDD.t86 VDD.t87 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X144 VDD.t85 VDD.t84 VDD.t85 VDD.t40 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X145 VSS.t139 VSS.t138 VSS.t139 VSS.t13 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X146 VSS.t137 VSS.t136 VSS.t137 VSS.t26 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X147 VSS.t135 VSS.t134 VSS.t135 VSS.t23 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X148 VDD.t83 VDD.t82 VDD.t83 VDD.t15 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X149 VDD.t81 VDD.t79 VDD.t81 VDD.t80 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X150 VDD.t78 VDD.t77 VDD.t78 VDD.t4 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X151 VSS.t133 VSS.t132 VSS.t133 VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X152 VSS.t131 VSS.t130 VSS.t131 VSS.t46 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X153 VDD a_n160_7781.t16 a_7622_1806# VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X154 VSS.t129 VSS.t128 VSS.t129 VSS.t41 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X155 VSS.t127 VSS.t126 VSS.t127 VSS.t38 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X156 VSS.t125 VSS.t124 VSS.t125 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X157 IBP a_5850_6555.t14 a_7656_7781# VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X158 VDD.t76 VDD.t74 VDD.t76 VDD.t75 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X159 a_13536_8547# IBP.t8 ITP.t1 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X160 a_13536_6615# IBP.t9 ITP.t2 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X161 a_7622_1806# a_n160_7781.t17 IBN.t0 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X162 VSS.t123 VSS.t122 VSS.t123 VSS.t29 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X163 VSS.t121 VSS.t120 VSS.t121 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X164 VSS.t119 VSS.t118 VSS.t119 VSS.t32 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X165 VSS.t117 VSS.t116 VSS.t117 VSS.t6 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X166 ITN a_12_588.t4 a_412_648# VSS.t18 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X167 VDD.t73 VDD.t72 VDD.t73 VDD.t7 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X168 VDD.t71 VDD.t70 VDD.t71 VDD.t40 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X169 a_7656_7781# a_5850_6555.t15 VSS.t2 VDD.t4 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X170 VDD.t69 VDD.t68 VDD.t69 VDD.t6 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X171 ITN IBN.t11 a_412_3730# VSS.t18 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X172 VSS.t115 VSS.t114 VSS.t115 VSS.t59 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X173 a_6250_9713# a_5850_6555.t16 VB.t1 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X174 VSS.t113 VSS.t112 VSS.t113 VSS.t26 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X175 VSS.t111 VSS.t110 VSS.t111 VSS.t21 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X176 VSS.t109 VSS.t108 VSS.t109 VSS.t23 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X177 VSS.t107 VSS.t106 VSS.t107 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X178 VSS.t105 VSS.t104 VSS.t105 VSS.t20 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X179 VSS.t103 VSS.t102 VSS.t103 VSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X180 VSS.t101 VSS.t100 VSS.t101 VSS.t49 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X181 VDD.t67 VDD.t66 VDD.t67 VDD.t6 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X182 VSS.t99 VSS.t98 VSS.t99 VSS.t7 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X183 a_12101_1806# a_11579_648.t19 a_5850_6555.t7 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X184 VDD.t65 VDD.t64 VDD.t65 VDD.t40 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X185 VSS.t97 VSS.t96 VSS.t97 VSS.t46 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X186 VSS.t95 VSS.t94 VSS.t95 VSS.t59 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X187 VDD.t63 VDD.t62 VDD.t63 VDD.t24 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X188 a_370_9713# a_n160_6615.t20 a_n160_7781.t6 VDD.t9 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X189 a_6250_8547# a_5850_6555.t18 IBP.t1 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X190 VSS.t93 VSS.t92 VSS.t93 VSS.t41 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X191 VSS.t91 VSS.t90 VSS.t91 VSS.t38 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X192 a_6250_6615# a_5850_6555.t19 VA.t1 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X193 a_13536_7781# a_12_588.t3 ITP.t5 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X194 ITN a_12_588.t2 a_412_2572# VSS.t18 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X195 VDD a_n160_6615.t21 a_370_9713# VDD.t10 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X196 VSS.t89 VSS.t88 VSS.t89 VSS.t13 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X197 VDD.t61 VDD.t60 VDD.t61 VDD.t21 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X198 a_12130_9713# IBP.t10 a_5850_6555.t0 VDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X199 VSS.t87 VSS.t86 VSS.t87 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X200 VSS a_5850_6555.t20 a_6250_8547# VDD.t2 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X201 VSS.t85 VSS.t84 VSS.t85 VSS.t49 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X202 VDD.t59 VDD.t58 VDD.t59 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X203 VSS.t83 VSS.t82 VSS.t83 VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X204 IBN a_n160_7781.t19 a_6218_2572# VSS.t5 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X205 VSS.t81 VSS.t80 VSS.t81 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X206 VDD.t57 VDD.t55 VDD.t57 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X207 VSS.t79 VSS.t78 VSS.t79 VSS.t29 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X208 VDD.t54 VDD.t52 VDD.t54 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X209 VSS.t77 VSS.t76 VSS.t77 VSS.t26 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X210 VSS.t75 VSS.t74 VSS.t75 VSS.t23 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X211 VSS.t73 VSS.t72 VSS.t73 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X212 VSS.t71 VSS.t70 VSS.t71 VSS.t6 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X213 a_370_8547# a_n160_6615.t2 a_n160_6615.t3 VDD.t9 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X214 a_370_6615# a_n160_6615.t4 a_n160_6615.t5 VDD.t9 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X215 VDD.t51 VDD.t50 VDD.t51 VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X216 VDD a_n160_6615.t22 a_370_8547# VDD.t10 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X217 VDD.t49 VDD.t48 VDD.t49 VDD.t21 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X218 VDD a_n160_6615.t23 a_370_6615# VDD.t10 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X219 a_12130_8547# a_12_588.t3 a_11579_648.t0 VDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X220 VSS.t69 VSS.t67 VSS.t69 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X221 VSS.t66 VSS.t65 VSS.t66 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X222 VDD.t47 VDD.t46 VDD.t47 VDD.t10 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X223 VDD.t45 VDD.t44 VDD.t45 VDD.t21 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X224 a_12130_6615# a_12_588.t3 a_11579_648.t0 VDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X225 VSS.t64 VSS.t63 VSS.t64 VSS.t32 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X226 VDD.t43 VDD.t42 VDD.t43 VDD.t2 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X227 a_7622_3730# a_n160_7781.t21 a_12_588.t2 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X228 VDD.t41 VDD.t39 VDD.t41 VDD.t40 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X229 VSS.t62 VSS.t61 VSS.t62 VSS.t49 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X230 a_6250_7781# a_5850_6555.t22 IBP.t2 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X231 VSS.t60 VSS.t58 VSS.t60 VSS.t59 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X232 VSS.t57 VSS.t56 VSS.t57 VSS.t32 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X233 VDD.t38 VDD.t36 VDD.t38 VDD.t37 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X234 VSS.t55 VSS.t54 VSS.t55 VSS.t18 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X235 VDD.t35 VDD.t34 VDD.t35 VDD.t9 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X236 VSS.t53 VSS.t51 VSS.t53 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X237 VSS a_5850_6555.t23 a_6250_7781# VDD.t2 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X238 a_1816_1806# a_12_588.t2 ITN.t4 VSS.t20 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X239 a_13505_1806# a_11579_648.t21 VSS.t11 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X240 VSS.t50 VSS.t48 VSS.t50 VSS.t49 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X241 VDD.t33 VDD.t32 VDD.t33 VDD.t10 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X242 VDD.t31 VDD.t30 VDD.t31 VDD.t21 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X243 VDD.t29 VDD.t28 VDD.t29 VDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X244 VDD.t27 VDD.t26 VDD.t27 VDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X245 VSS.t47 VSS.t45 VSS.t47 VSS.t46 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X246 VSS.t44 VSS.t43 VSS.t44 VSS.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X247 VSS.t42 VSS.t40 VSS.t42 VSS.t41 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X248 VSS.t39 VSS.t37 VSS.t39 VSS.t38 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X249 a_12101_3730# a_11579_648.t22 a_5850_6555.t5 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X250 VDD a_n160_7781.t22 a_7622_2572# VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X251 a_7622_2572# a_n160_7781.t23 IBN.t1 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X252 a_370_7781# a_n160_6615.t24 a_n160_7781.t7 VDD.t9 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X253 VDD.t25 VDD.t23 VDD.t25 VDD.t24 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X254 VSS a_11579_648.t23 a_12101_648# VSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X255 VSS.t36 VSS.t34 VSS.t36 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X256 VDD a_n160_6615.t25 a_370_7781# VDD.t10 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X257 VSS.t33 VSS.t31 VSS.t33 VSS.t32 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X258 VDD.t22 VDD.t20 VDD.t22 VDD.t21 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X259 VDD.t19 VDD.t18 VDD.t19 VDD.t4 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X260 a_12130_7781# IBP.t11 a_5850_6555.t3 VDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X261 VSS a_11579_648.t24 a_12101_1806# VSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X262 a_412_648# a_12_588.t4 a_n160_6615.t11 VSS.t19 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X263 VSS.t30 VSS.t28 VSS.t30 VSS.t29 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X264 VSS.t27 VSS.t25 VSS.t27 VSS.t26 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X265 VSS.t24 VSS.t22 VSS.t24 VSS.t23 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
R0 IBP.n21 IBP.n20 9.90372
R1 IBP.n14 IBP.t8 8.44198
R2 IBP.n14 IBP.t6 8.44198
R3 IBP.n2 IBP.t9 8.44198
R4 IBP.n2 IBP.t7 8.44198
R5 IBP.n13 IBP.t10 8.10925
R6 IBP.n5 IBP.t11 8.10925
R7 IBP.n18 IBP.t4 8.10567
R8 IBP.n8 IBP.t5 8.10567
R9 IBP.n22 IBP.n1 4.84877
R10 IBP.n19 IBP.n18 4.63432
R11 IBP.n9 IBP.n8 4.63432
R12 IBP.n1 IBP.t1 3.65383
R13 IBP.n23 IBP.n0 3.65146
R14 IBP.n1 IBP.t2 3.57094
R15 IBP IBP.n24 3.4916
R16 IBP.n20 IBP.n19 3.37487
R17 IBP.n10 IBP.n9 3.37487
R18 IBP.n22 IBP.n21 3.11372
R19 IBP.n3 IBP.n2 2.86385
R20 IBP.n15 IBP.n14 2.85082
R21 IBP.n23 IBP.n22 2.71171
R22 IBP.n17 IBP.n16 2.3531
R23 IBP.n7 IBP.n6 2.34007
R24 IBP.n10 IBP.n3 2.30075
R25 IBP.n16 IBP.n13 2.28392
R26 IBP.n6 IBP.n5 2.2709
R27 IBP.n17 IBP.n12 2.25205
R28 IBP.n7 IBP.n4 2.25205
R29 IBP.n15 IBP.n11 2.2505
R30 IBP.n13 IBP.n12 2.09285
R31 IBP.n5 IBP.n4 2.09285
R32 IBP.n16 IBP.n15 1.28862
R33 IBP.n6 IBP.n3 1.28862
R34 IBP.n11 IBP.n10 0.670625
R35 IBP.n21 IBP 0.372239
R36 IBP.n19 IBP.n12 0.234207
R37 IBP.n9 IBP.n4 0.234207
R38 IBP IBP.n23 0.0822105
R39 IBP.n20 IBP.n11 0.054875
R40 IBP.n18 IBP.n17 0.00997368
R41 IBP.n8 IBP.n7 0.00997368
R42 ITP.n9 ITP.t7 6.54387
R43 ITP.n1 ITP.t2 6.39955
R44 ITP.n1 ITP.n0 5.83655
R45 ITP.n7 ITP.n1 4.03827
R46 ITP.n5 ITP.n3 3.73554
R47 ITP.n2 ITP.t1 3.73554
R48 ITP.n5 ITP.n4 3.57923
R49 ITP.n2 ITP.t5 3.57923
R50 ITP ITP.n10 3.48212
R51 ITP.n7 ITP.n6 3.45552
R52 ITP.n9 ITP.n8 3.35988
R53 ITP.n6 ITP.n2 2.58435
R54 ITP ITP.n9 2.51007
R55 ITP.n6 ITP.n5 2.22754
R56 ITP.n8 ITP.n7 0.780125
R57 ITP.n8 ITP 0.4175
R58 VDD.n178 VDD.n21 477.971
R59 VDD.n88 VDD.n46 477.971
R60 VDD.n217 VDD.n10 477.971
R61 VDD.n175 VDD.n5 470.842
R62 VDD.n83 VDD.n27 470.842
R63 VDD.n213 VDD.n9 470.842
R64 VDD.n178 VDD.n5 470.842
R65 VDD.n88 VDD.n27 470.842
R66 VDD.n213 VDD.n10 470.842
R67 VDD.n175 VDD.n21 469.683
R68 VDD.n83 VDD.n46 469.683
R69 VDD.n217 VDD.n9 469.683
R70 VDD.t7 VDD.t123 142.93
R71 VDD.t5 VDD.t53 142.93
R72 VDD.t80 VDD.t3 142.93
R73 VDD.t1 VDD.t100 142.93
R74 VDD.t21 VDD.t149 142.93
R75 VDD.t9 VDD.t93 142.93
R76 VDD.t123 VDD.t40 96.8792
R77 VDD.t6 VDD.t7 96.8792
R78 VDD.t8 VDD.t5 96.8792
R79 VDD.t53 VDD.t142 96.8792
R80 VDD.t75 VDD.t80 96.8792
R81 VDD.t3 VDD.t4 96.8792
R82 VDD.t2 VDD.t1 96.8792
R83 VDD.t100 VDD.t24 96.8792
R84 VDD.t56 VDD.t21 96.8792
R85 VDD.t149 VDD.t15 96.8792
R86 VDD.t10 VDD.t9 96.8792
R87 VDD.t93 VDD.t37 96.8792
R88 VDD.t40 VDD.n46 81.1238
R89 VDD.t37 VDD.n213 81.1238
R90 VDD.t142 VDD.n86 81.017
R91 VDD.n85 VDD.t75 81.017
R92 VDD.t24 VDD.n11 81.017
R93 VDD.n216 VDD.t56 81.017
R94 VDD.n84 VDD.t6 70.2717
R95 VDD.n176 VDD.t4 70.2717
R96 VDD.t15 VDD.n215 70.2717
R97 VDD.n87 VDD.t8 64.1315
R98 VDD.n177 VDD.t2 64.1315
R99 VDD.n214 VDD.t10 64.1315
R100 VDD.n86 VDD.n85 24.5613
R101 VDD.n216 VDD.n11 24.5613
R102 VDD.n87 VDD.n84 8.52856
R103 VDD.n177 VDD.n176 8.52856
R104 VDD.n215 VDD.n214 8.52856
R105 VDD.n225 VDD.t211 8.10567
R106 VDD.n225 VDD.t55 8.10567
R107 VDD.n222 VDD.t60 8.10567
R108 VDD.n222 VDD.t221 8.10567
R109 VDD.n221 VDD.t48 8.10567
R110 VDD.n221 VDD.t209 8.10567
R111 VDD.n185 VDD.t20 8.10567
R112 VDD.n185 VDD.t163 8.10567
R113 VDD.n186 VDD.t44 8.10567
R114 VDD.n186 VDD.t205 8.10567
R115 VDD.n190 VDD.t30 8.10567
R116 VDD.n190 VDD.t183 8.10567
R117 VDD.n225 VDD.t62 8.10567
R118 VDD.n225 VDD.t125 8.10567
R119 VDD.n222 VDD.t23 8.10567
R120 VDD.n222 VDD.t169 8.10567
R121 VDD.n221 VDD.t217 8.10567
R122 VDD.n221 VDD.t144 8.10567
R123 VDD.n185 VDD.t179 8.10567
R124 VDD.n185 VDD.t99 8.10567
R125 VDD.n186 VDD.t215 8.10567
R126 VDD.n186 VDD.t137 8.10567
R127 VDD.n190 VDD.t197 8.10567
R128 VDD.n190 VDD.t112 8.10567
R129 VDD.n170 VDD.t159 8.10567
R130 VDD.n121 VDD.t189 8.10567
R131 VDD.n22 VDD.t18 8.10567
R132 VDD.n117 VDD.t58 8.10567
R133 VDD.n125 VDD.t102 8.10567
R134 VDD.n123 VDD.t46 8.10567
R135 VDD.n164 VDD.t82 8.10567
R136 VDD.n122 VDD.t148 8.10567
R137 VDD.n132 VDD.t36 8.10567
R138 VDD.n132 VDD.t207 8.10567
R139 VDD.n130 VDD.t161 8.10567
R140 VDD.n130 VDD.t165 8.10567
R141 VDD.n129 VDD.t135 8.10567
R142 VDD.n129 VDD.t139 8.10567
R143 VDD.n210 VDD.t90 8.10567
R144 VDD.n210 VDD.t92 8.10567
R145 VDD.n209 VDD.t129 8.10567
R146 VDD.n209 VDD.t133 8.10567
R147 VDD.n207 VDD.t108 8.10567
R148 VDD.n207 VDD.t110 8.10567
R149 VDD.n78 VDD.t28 8.10567
R150 VDD.n77 VDD.t104 8.10567
R151 VDD.n47 VDD.t68 8.10567
R152 VDD.n73 VDD.t120 8.10567
R153 VDD.n70 VDD.t191 8.10567
R154 VDD.n70 VDD.t39 8.10567
R155 VDD.n68 VDD.t199 8.10567
R156 VDD.n68 VDD.t114 8.10567
R157 VDD.n67 VDD.t175 8.10567
R158 VDD.n67 VDD.t88 8.10567
R159 VDD.n63 VDD.t122 8.10567
R160 VDD.n63 VDD.t64 8.10567
R161 VDD.n62 VDD.t173 8.10567
R162 VDD.n62 VDD.t84 8.10567
R163 VDD.n60 VDD.t151 8.10567
R164 VDD.n60 VDD.t70 8.10567
R165 VDD.n44 VDD.t26 8.10567
R166 VDD.n91 VDD.t187 8.10567
R167 VDD.n55 VDD.t66 8.10567
R168 VDD.n54 VDD.t72 8.10567
R169 VDD.n19 VDD.t50 8.10567
R170 VDD.n181 VDD.t42 8.10567
R171 VDD.n32 VDD.t77 8.10567
R172 VDD.n35 VDD.t97 8.10567
R173 VDD.n112 VDD.t79 8.10567
R174 VDD.n112 VDD.t177 8.10567
R175 VDD.n109 VDD.t219 8.10567
R176 VDD.n109 VDD.t146 8.10567
R177 VDD.n108 VDD.t203 8.10567
R178 VDD.n108 VDD.t118 8.10567
R179 VDD.n102 VDD.t157 8.10567
R180 VDD.n102 VDD.t74 8.10567
R181 VDD.n101 VDD.t201 8.10567
R182 VDD.n101 VDD.t116 8.10567
R183 VDD.n98 VDD.t181 8.10567
R184 VDD.n98 VDD.t95 8.10567
R185 VDD.n112 VDD.t141 8.10567
R186 VDD.n112 VDD.t52 8.10567
R187 VDD.n109 VDD.t213 8.10567
R188 VDD.n109 VDD.t155 8.10567
R189 VDD.n108 VDD.t195 8.10567
R190 VDD.n108 VDD.t131 8.10567
R191 VDD.n102 VDD.t153 8.10567
R192 VDD.n102 VDD.t86 8.10567
R193 VDD.n101 VDD.t193 8.10567
R194 VDD.n101 VDD.t127 8.10567
R195 VDD.n98 VDD.t167 8.10567
R196 VDD.n98 VDD.t106 8.10567
R197 VDD.n17 VDD.t34 8.10567
R198 VDD.n202 VDD.t32 8.10567
R199 VDD.n18 VDD.t171 8.10567
R200 VDD.n196 VDD.t185 8.10567
R201 VDD.n42 VDD.n41 5.76894
R202 VDD.n41 VDD.n40 5.33948
R203 VDD.n154 VDD.n153 4.61205
R204 VDD.n143 VDD.n142 4.61205
R205 VDD.n42 VDD.n36 4.57315
R206 VDD.n43 VDD.n42 4.56231
R207 VDD.n147 VDD.n145 4.5005
R208 VDD.n140 VDD.n138 4.5005
R209 VDD.n158 VDD.n157 4.5005
R210 VDD.n157 VDD.n126 4.5005
R211 VDD.n136 VDD.n124 4.5005
R212 VDD.n136 VDD.n135 4.5005
R213 VDD.n137 VDD.t17 4.00848
R214 VDD.n142 VDD.n141 4.00554
R215 VDD.n40 VDD.t225 3.8555
R216 VDD.n39 VDD.n37 3.85313
R217 VDD.n137 VDD.t227 3.78097
R218 VDD.n148 VDD.t224 3.78097
R219 VDD.n147 VDD.n146 3.77818
R220 VDD.n140 VDD.n139 3.77818
R221 VDD.n39 VDD.n38 3.68497
R222 VDD.n40 VDD.t226 3.68261
R223 VDD.n144 VDD.n143 3.54958
R224 VDD.n150 VDD.n144 3.27995
R225 VDD.n169 VDD.t160 3.20383
R226 VDD.n173 VDD.t190 3.20383
R227 VDD.n120 VDD.t19 3.20383
R228 VDD.n116 VDD.t59 3.20383
R229 VDD.n134 VDD.t103 3.20383
R230 VDD.n161 VDD.t47 3.20383
R231 VDD.n163 VDD.t83 3.20383
R232 VDD.n167 VDD.t150 3.20383
R233 VDD.n149 VDD.t16 3.20383
R234 VDD.n152 VDD.n151 3.20383
R235 VDD.t29 VDD.n23 3.20383
R236 VDD.n81 VDD.t105 3.20383
R237 VDD.n76 VDD.t69 3.20383
R238 VDD.n72 VDD.t121 3.20383
R239 VDD.n94 VDD.t27 3.20383
R240 VDD.n90 VDD.t188 3.20383
R241 VDD.t67 VDD.n45 3.20383
R242 VDD.n58 VDD.t73 3.20383
R243 VDD.n184 VDD.t51 3.20383
R244 VDD.n180 VDD.t43 3.20383
R245 VDD.t78 VDD.n20 3.20383
R246 VDD.t98 VDD.n31 3.20383
R247 VDD.n205 VDD.t35 3.20383
R248 VDD.n201 VDD.t33 3.20383
R249 VDD.n199 VDD.t172 3.20383
R250 VDD.n195 VDD.t186 3.20383
R251 VDD.n155 VDD.n154 3.2012
R252 VDD.n150 VDD.n149 3.1154
R253 VDD.n148 VDD.n145 2.65924
R254 VDD.n138 VDD.n137 2.65924
R255 VDD.n152 VDD.n150 2.61766
R256 VDD.n34 VDD.n33 1.73383
R257 VDD.n183 VDD.n182 1.73383
R258 VDD.n57 VDD.n56 1.73383
R259 VDD.n93 VDD.n92 1.73383
R260 VDD.n75 VDD.n74 1.73383
R261 VDD.n80 VDD.n79 1.73383
R262 VDD.n198 VDD.n197 1.73383
R263 VDD.n204 VDD.n203 1.73383
R264 VDD.n166 VDD.n165 1.73383
R265 VDD.n160 VDD.n159 1.73383
R266 VDD.n119 VDD.n118 1.73383
R267 VDD.n172 VDD.n171 1.73383
R268 VDD.n156 VDD.n155 1.59478
R269 VDD.n41 VDD.n39 1.49396
R270 VDD.t190 VDD.n172 1.4705
R271 VDD.n172 VDD.t160 1.4705
R272 VDD.n119 VDD.t59 1.4705
R273 VDD.t19 VDD.n119 1.4705
R274 VDD.t47 VDD.n160 1.4705
R275 VDD.n160 VDD.t103 1.4705
R276 VDD.t150 VDD.n166 1.4705
R277 VDD.n166 VDD.t83 1.4705
R278 VDD.t105 VDD.n80 1.4705
R279 VDD.n80 VDD.t29 1.4705
R280 VDD.n75 VDD.t121 1.4705
R281 VDD.t69 VDD.n75 1.4705
R282 VDD.n93 VDD.t188 1.4705
R283 VDD.t27 VDD.n93 1.4705
R284 VDD.t73 VDD.n57 1.4705
R285 VDD.n57 VDD.t67 1.4705
R286 VDD.n183 VDD.t43 1.4705
R287 VDD.t51 VDD.n183 1.4705
R288 VDD.n33 VDD.t98 1.4705
R289 VDD.n33 VDD.t78 1.4705
R290 VDD.n204 VDD.t33 1.4705
R291 VDD.t35 VDD.n204 1.4705
R292 VDD.n198 VDD.t186 1.4705
R293 VDD.t172 VDD.n198 1.4705
R294 VDD.n0 VDD.t57 1.00929
R295 VDD.n3 VDD.t222 1.00929
R296 VDD.n4 VDD.t210 1.00929
R297 VDD.n6 VDD.t164 1.00929
R298 VDD.n187 VDD.t206 1.00929
R299 VDD.n191 VDD.t184 1.00929
R300 VDD.n1 VDD.t126 1.00929
R301 VDD.n223 VDD.t170 1.00929
R302 VDD.n219 VDD.t145 1.00929
R303 VDD.n7 VDD.t101 1.00929
R304 VDD.n188 VDD.t138 1.00929
R305 VDD.n192 VDD.t113 1.00929
R306 VDD.n127 VDD.t208 1.00929
R307 VDD.n128 VDD.t166 1.00929
R308 VDD.n12 VDD.t140 1.00929
R309 VDD.n14 VDD.t94 1.00929
R310 VDD.n15 VDD.t134 1.00929
R311 VDD.n16 VDD.t111 1.00929
R312 VDD.n48 VDD.t41 1.00929
R313 VDD.n49 VDD.t115 1.00929
R314 VDD.n50 VDD.t89 1.00929
R315 VDD.n51 VDD.t65 1.00929
R316 VDD.n52 VDD.t85 1.00929
R317 VDD.n53 VDD.t71 1.00929
R318 VDD.n24 VDD.t178 1.00929
R319 VDD.n25 VDD.t147 1.00929
R320 VDD.n26 VDD.t119 1.00929
R321 VDD.n28 VDD.t76 1.00929
R322 VDD.n29 VDD.t117 1.00929
R323 VDD.n30 VDD.t96 1.00929
R324 VDD.n113 VDD.t54 1.00929
R325 VDD.n110 VDD.t156 1.00929
R326 VDD.n106 VDD.t132 1.00929
R327 VDD.n103 VDD.t87 1.00929
R328 VDD.n99 VDD.t128 1.00929
R329 VDD.n96 VDD.t107 1.00929
R330 VDD.n0 VDD.t212 1.00871
R331 VDD.n3 VDD.t61 1.00871
R332 VDD.n4 VDD.t49 1.00871
R333 VDD.n6 VDD.t22 1.00871
R334 VDD.n187 VDD.t45 1.00871
R335 VDD.n191 VDD.t31 1.00871
R336 VDD.n1 VDD.t63 1.00871
R337 VDD.n223 VDD.t25 1.00871
R338 VDD.n219 VDD.t218 1.00871
R339 VDD.n7 VDD.t180 1.00871
R340 VDD.n188 VDD.t216 1.00871
R341 VDD.n192 VDD.t198 1.00871
R342 VDD.n127 VDD.t38 1.00871
R343 VDD.n128 VDD.t162 1.00871
R344 VDD.n12 VDD.t136 1.00871
R345 VDD.n14 VDD.t91 1.00871
R346 VDD.n15 VDD.t130 1.00871
R347 VDD.n16 VDD.t109 1.00871
R348 VDD.n48 VDD.t192 1.00871
R349 VDD.n49 VDD.t200 1.00871
R350 VDD.n50 VDD.t176 1.00871
R351 VDD.n51 VDD.t124 1.00871
R352 VDD.n52 VDD.t174 1.00871
R353 VDD.n53 VDD.t152 1.00871
R354 VDD.n24 VDD.t81 1.00871
R355 VDD.n25 VDD.t220 1.00871
R356 VDD.n26 VDD.t204 1.00871
R357 VDD.n28 VDD.t158 1.00871
R358 VDD.n29 VDD.t202 1.00871
R359 VDD.n30 VDD.t182 1.00871
R360 VDD.n113 VDD.t143 1.00871
R361 VDD.n110 VDD.t214 1.00871
R362 VDD.n106 VDD.t196 1.00871
R363 VDD.n103 VDD.t154 1.00871
R364 VDD.n99 VDD.t194 1.00871
R365 VDD.n96 VDD.t168 1.00871
R366 VDD.n149 VDD.n148 0.805146
R367 VDD.n153 VDD.n152 0.80221
R368 VDD.n97 VDD.n96 0.468749
R369 VDD.n100 VDD.n99 0.468749
R370 VDD.n104 VDD.n103 0.468749
R371 VDD.n107 VDD.n106 0.468749
R372 VDD.n111 VDD.n110 0.468749
R373 VDD.n114 VDD.n113 0.468749
R374 VDD.n97 VDD.n30 0.468749
R375 VDD.n100 VDD.n29 0.468749
R376 VDD.n104 VDD.n28 0.468749
R377 VDD.n107 VDD.n26 0.468749
R378 VDD.n111 VDD.n25 0.468749
R379 VDD.n114 VDD.n24 0.468749
R380 VDD.n59 VDD.n53 0.468749
R381 VDD.n61 VDD.n52 0.468749
R382 VDD.n64 VDD.n51 0.468749
R383 VDD.n66 VDD.n50 0.468749
R384 VDD.n69 VDD.n49 0.468749
R385 VDD.n71 VDD.n48 0.468749
R386 VDD.n206 VDD.n16 0.468749
R387 VDD.n208 VDD.n15 0.468749
R388 VDD.n211 VDD.n14 0.468749
R389 VDD.n13 VDD.n12 0.468749
R390 VDD.n131 VDD.n128 0.468749
R391 VDD.n133 VDD.n127 0.468749
R392 VDD.n193 VDD.n192 0.468749
R393 VDD.n189 VDD.n188 0.468749
R394 VDD.n8 VDD.n7 0.468749
R395 VDD.n220 VDD.n219 0.468749
R396 VDD.n224 VDD.n223 0.468749
R397 VDD.n2 VDD.n1 0.468749
R398 VDD.n193 VDD.n191 0.468749
R399 VDD.n189 VDD.n187 0.468749
R400 VDD.n8 VDD.n6 0.468749
R401 VDD.n220 VDD.n4 0.468749
R402 VDD.n224 VDD.n3 0.468749
R403 VDD.n2 VDD.n0 0.468749
R404 VDD.n155 VDD.n144 0.3755
R405 VDD.n154 VDD.n145 0.157683
R406 VDD.n143 VDD.n138 0.157683
R407 VDD.n83 VDD.n82 0.10728
R408 VDD.n84 VDD.n83 0.10728
R409 VDD.n65 VDD.n46 0.10728
R410 VDD.n105 VDD.n27 0.10728
R411 VDD.n86 VDD.n27 0.10728
R412 VDD.n105 VDD.n21 0.10728
R413 VDD.n85 VDD.n21 0.10728
R414 VDD.n213 VDD.n212 0.10728
R415 VDD.n162 VDD.n9 0.10728
R416 VDD.n215 VDD.n9 0.10728
R417 VDD.n175 VDD.n174 0.10728
R418 VDD.n176 VDD.n175 0.10728
R419 VDD.n218 VDD.n5 0.10728
R420 VDD.n11 VDD.n5 0.10728
R421 VDD.n218 VDD.n217 0.10728
R422 VDD.n217 VDD.n216 0.10728
R423 VDD.n89 VDD.n88 0.1055
R424 VDD.n88 VDD.n87 0.1055
R425 VDD.n179 VDD.n178 0.1055
R426 VDD.n178 VDD.n177 0.1055
R427 VDD.n200 VDD.n10 0.1055
R428 VDD.n214 VDD.n10 0.1055
R429 VDD.n70 VDD.n69 0.0382419
R430 VDD.n61 VDD.n60 0.0382419
R431 VDD.n132 VDD.n131 0.0382419
R432 VDD.n208 VDD.n207 0.0382419
R433 VDD.n68 VDD.n67 0.0364748
R434 VDD.n63 VDD.n62 0.0364748
R435 VDD.n130 VDD.n129 0.0364748
R436 VDD.n210 VDD.n209 0.0364748
R437 VDD.n73 VDD.n72 0.0346711
R438 VDD.n74 VDD.n73 0.0346711
R439 VDD.n74 VDD.n47 0.0346711
R440 VDD.n76 VDD.n47 0.0346711
R441 VDD.n81 VDD.n77 0.0346711
R442 VDD.n79 VDD.n77 0.0346711
R443 VDD.n79 VDD.n78 0.0346711
R444 VDD.n78 VDD.n23 0.0346711
R445 VDD.n167 VDD.n122 0.0346711
R446 VDD.n165 VDD.n122 0.0346711
R447 VDD.n165 VDD.n164 0.0346711
R448 VDD.n164 VDD.n163 0.0346711
R449 VDD.n161 VDD.n123 0.0346711
R450 VDD.n159 VDD.n123 0.0346711
R451 VDD.n117 VDD.n116 0.0346711
R452 VDD.n118 VDD.n117 0.0346711
R453 VDD.n118 VDD.n22 0.0346711
R454 VDD.n120 VDD.n22 0.0346711
R455 VDD.n173 VDD.n121 0.0346711
R456 VDD.n171 VDD.n121 0.0346711
R457 VDD.n171 VDD.n170 0.0346711
R458 VDD.n170 VDD.n169 0.0346711
R459 VDD.n59 VDD.n58 0.0308563
R460 VDD.n206 VDD.n205 0.0308563
R461 VDD.n72 VDD.n71 0.0308128
R462 VDD.n134 VDD.n133 0.0308128
R463 VDD.n159 VDD.n158 0.0302193
R464 VDD.n35 VDD.n34 0.0293162
R465 VDD.n34 VDD.n32 0.0293162
R466 VDD.n32 VDD.n20 0.0293162
R467 VDD.n181 VDD.n180 0.0293162
R468 VDD.n182 VDD.n181 0.0293162
R469 VDD.n182 VDD.n19 0.0293162
R470 VDD.n184 VDD.n19 0.0293162
R471 VDD.n58 VDD.n54 0.0293162
R472 VDD.n56 VDD.n54 0.0293162
R473 VDD.n56 VDD.n55 0.0293162
R474 VDD.n55 VDD.n45 0.0293162
R475 VDD.n91 VDD.n90 0.0293162
R476 VDD.n92 VDD.n91 0.0293162
R477 VDD.n92 VDD.n44 0.0293162
R478 VDD.n94 VDD.n44 0.0293162
R479 VDD.n196 VDD.n195 0.0293162
R480 VDD.n197 VDD.n196 0.0293162
R481 VDD.n197 VDD.n18 0.0293162
R482 VDD.n199 VDD.n18 0.0293162
R483 VDD.n202 VDD.n201 0.0293162
R484 VDD.n203 VDD.n202 0.0293162
R485 VDD.n203 VDD.n17 0.0293162
R486 VDD.n205 VDD.n17 0.0293162
R487 VDD.n115 VDD.n23 0.0284144
R488 VDD.n168 VDD.n167 0.0284144
R489 VDD.n116 VDD.n115 0.0284144
R490 VDD.n169 VDD.n168 0.0284144
R491 VDD.n156 VDD.n136 0.0271036
R492 VDD.n66 VDD.n65 0.0270708
R493 VDD.n212 VDD.n13 0.0270708
R494 VDD.n135 VDD.n134 0.0240829
R495 VDD.n194 VDD.n184 0.02404
R496 VDD.n95 VDD.n94 0.02404
R497 VDD.n195 VDD.n194 0.02404
R498 VDD.n36 VDD.n35 0.0232283
R499 VDD.n65 VDD.n64 0.0222742
R500 VDD.n212 VDD.n211 0.0222742
R501 VDD.n157 VDD.n156 0.0199738
R502 VDD.n71 VDD.n70 0.0193079
R503 VDD.n69 VDD.n68 0.0193079
R504 VDD.n67 VDD.n66 0.0193079
R505 VDD.n64 VDD.n63 0.0193079
R506 VDD.n62 VDD.n61 0.0193079
R507 VDD.n60 VDD.n59 0.0193079
R508 VDD.n133 VDD.n132 0.0193079
R509 VDD.n131 VDD.n130 0.0193079
R510 VDD.n129 VDD.n13 0.0193079
R511 VDD.n211 VDD.n210 0.0193079
R512 VDD.n209 VDD.n208 0.0193079
R513 VDD.n207 VDD.n206 0.0193079
R514 VDD.n112 VDD.n111 0.0192265
R515 VDD.n100 VDD.n98 0.0192265
R516 VDD.n225 VDD.n224 0.0192265
R517 VDD.n190 VDD.n189 0.0192265
R518 VDD.n179 VDD.n20 0.0185609
R519 VDD.n89 VDD.n45 0.0185609
R520 VDD.n200 VDD.n199 0.0185609
R521 VDD.n109 VDD.n108 0.0183497
R522 VDD.n102 VDD.n101 0.0183497
R523 VDD.n222 VDD.n221 0.0183497
R524 VDD.n186 VDD.n185 0.0183497
R525 VDD.n82 VDD.n81 0.0175856
R526 VDD.n162 VDD.n161 0.0175856
R527 VDD.n174 VDD.n173 0.0175856
R528 VDD.n95 VDD.n43 0.0175462
R529 VDD.n82 VDD.n76 0.0159011
R530 VDD.n163 VDD.n162 0.0159011
R531 VDD.n174 VDD.n120 0.0159011
R532 VDD.n107 VDD.n105 0.0136837
R533 VDD.n220 VDD.n218 0.0136837
R534 VDD.n105 VDD.n104 0.0113038
R535 VDD.n218 VDD.n8 0.0113038
R536 VDD.n126 VDD.n125 0.0109679
R537 VDD.n180 VDD.n179 0.00983484
R538 VDD.n90 VDD.n89 0.00983484
R539 VDD.n201 VDD.n200 0.00983484
R540 VDD.n114 VDD.n112 0.00983194
R541 VDD.n111 VDD.n109 0.00983194
R542 VDD.n108 VDD.n107 0.00983194
R543 VDD.n104 VDD.n102 0.00983194
R544 VDD.n101 VDD.n100 0.00983194
R545 VDD.n98 VDD.n97 0.00983194
R546 VDD.n224 VDD.n222 0.00983194
R547 VDD.n221 VDD.n220 0.00983194
R548 VDD.n185 VDD.n8 0.00983194
R549 VDD.n189 VDD.n186 0.00983194
R550 VDD.n193 VDD.n190 0.00983194
R551 VDD VDD.n225 0.00760856
R552 VDD.n43 VDD.n31 0.0069938
R553 VDD.n36 VDD.n31 0.00658794
R554 VDD.n153 VDD.n147 0.00523684
R555 VDD.n142 VDD.n140 0.00523684
R556 VDD.n125 VDD.n124 0.00483155
R557 VDD.n97 VDD.n95 0.00388205
R558 VDD.n194 VDD.n193 0.00388205
R559 VDD VDD.n2 0.00272338
R560 VDD.n115 VDD.n114 0.00168998
R561 VDD.n168 VDD.n2 0.00168998
R562 VDD.n158 VDD.n124 0.000620321
R563 VDD.n135 VDD.n126 0.000620321
R564 IBN.n23 IBN.n22 9.58265
R565 IBN.n1 IBN.t8 8.41259
R566 IBN.n12 IBN.t6 8.41259
R567 IBN.n1 IBN.t7 8.3889
R568 IBN.n12 IBN.t5 8.3889
R569 IBN.n3 IBN.t11 8.06917
R570 IBN.n2 IBN.t9 8.06917
R571 IBN.n15 IBN.t10 8.06917
R572 IBN.n13 IBN.t4 8.06917
R573 IBN.n4 IBN.n3 4.64616
R574 IBN.n16 IBN.n15 4.64616
R575 IBN.n7 IBN.n0 4.64379
R576 IBN.n19 IBN.n14 4.64379
R577 IBN.n6 IBN.n5 4.5005
R578 IBN.n18 IBN.n17 4.5005
R579 IBN.n28 IBN.t0 3.84484
R580 IBN.n26 IBN.n25 3.84484
R581 IBN.n26 IBN.n24 3.69326
R582 IBN IBN.t1 3.64116
R583 IBN.n27 IBN.n23 3.62732
R584 IBN.n10 IBN.n0 3.48328
R585 IBN.n14 IBN.n11 3.43191
R586 IBN.n9 IBN.n1 2.79852
R587 IBN.n21 IBN.n12 2.79497
R588 IBN.n20 IBN.n19 2.34718
R589 IBN.n8 IBN.n7 2.34362
R590 IBN.n20 IBN.n13 2.27585
R591 IBN.n8 IBN.n2 2.2723
R592 IBN.n22 IBN.n21 2.2505
R593 IBN.n10 IBN.n9 2.2505
R594 IBN.n4 IBN.n2 2.01635
R595 IBN.n16 IBN.n13 2.01635
R596 IBN.n9 IBN.n8 1.34566
R597 IBN.n21 IBN.n20 1.34566
R598 IBN.n11 IBN.n10 0.671
R599 IBN.n23 IBN 0.343707
R600 IBN.n27 IBN.n26 0.188652
R601 IBN.n5 IBN.n0 0.157683
R602 IBN.n5 IBN.n4 0.157683
R603 IBN.n17 IBN.n14 0.157683
R604 IBN.n17 IBN.n16 0.157683
R605 IBN.n28 IBN.n27 0.132718
R606 IBN.n22 IBN.n11 0.053
R607 IBN IBN.n28 0.0526053
R608 IBN.n7 IBN.n6 0.00405263
R609 IBN.n19 IBN.n18 0.00405263
R610 IBN.n6 IBN.n3 0.00168421
R611 IBN.n18 IBN.n15 0.00168421
R612 a_n160_7781.n2 a_n160_7781.t9 12.8637
R613 a_n160_7781.n1 a_n160_7781.t6 10.7018
R614 a_n160_7781.n1 a_n160_7781.t1 10.1659
R615 a_n160_7781.n1 a_n160_7781.n3 9.64387
R616 a_n160_7781.n1 a_n160_7781.n5 9.27665
R617 a_n160_7781.n1 a_n160_7781.n2 8.75198
R618 a_n160_7781.n2 a_n160_7781.t10 8.14051
R619 a_n160_7781.n2 a_n160_7781.t15 8.14051
R620 a_n160_7781.n2 a_n160_7781.t8 8.14051
R621 a_n160_7781.n2 a_n160_7781.t14 8.14051
R622 a_n160_7781.n2 a_n160_7781.t21 8.06917
R623 a_n160_7781.n2 a_n160_7781.t23 8.06917
R624 a_n160_7781.n2 a_n160_7781.t19 8.06917
R625 a_n160_7781.n2 a_n160_7781.t18 8.06917
R626 a_n160_7781.n2 a_n160_7781.t17 8.06917
R627 a_n160_7781.n2 a_n160_7781.t13 8.06917
R628 a_n160_7781.n2 a_n160_7781.t12 8.06917
R629 a_n160_7781.n0 a_n160_7781.t3 7.94068
R630 a_n160_7781.n1 a_n160_7781.t7 7.72524
R631 a_n160_7781.n0 a_n160_7781.n4 7.22855
R632 a_n160_7781.n6 a_n160_7781.n1 7.17942
R633 a_n160_7781.t22 a_n160_7781.n2 8.33649
R634 a_n160_7781.n2 a_n160_7781.t20 8.33649
R635 a_n160_7781.t11 a_n160_7781.n2 8.33556
R636 a_n160_7781.n2 a_n160_7781.t16 8.33556
R637 a_n160_7781.n1 a_n160_7781.n0 7.46075
R638 VSS.n153 VSS.n14 523.342
R639 VSS.n104 VSS.n20 523.342
R640 VSS.n206 VSS.n8 523.342
R641 VSS.n147 VSS.n15 521.869
R642 VSS.n107 VSS.n38 521.869
R643 VSS.n209 VSS.n7 521.869
R644 VSS.n147 VSS.n14 519.659
R645 VSS.n104 VSS.n38 519.659
R646 VSS.n206 VSS.n7 519.659
R647 VSS.n153 VSS.n15 516.342
R648 VSS.n107 VSS.n20 516.342
R649 VSS.n209 VSS.n8 516.342
R650 VSS.t0 VSS.t38 407.8
R651 VSS.t1 VSS.t52 407.8
R652 VSS.t4 VSS.t32 407.8
R653 VSS.t35 VSS.t6 407.8
R654 VSS.t41 VSS.t21 407.8
R655 VSS.t19 VSS.t68 407.8
R656 VSS.t38 VSS.t23 277.82
R657 VSS.t7 VSS.t0 277.82
R658 VSS.t13 VSS.t1 277.82
R659 VSS.t52 VSS.t49 277.82
R660 VSS.t32 VSS.t46 277.82
R661 VSS.t3 VSS.t4 277.82
R662 VSS.t6 VSS.t5 277.82
R663 VSS.t29 VSS.t35 277.82
R664 VSS.t26 VSS.t41 277.82
R665 VSS.t21 VSS.t20 277.82
R666 VSS.t18 VSS.t19 277.82
R667 VSS.t68 VSS.t59 277.82
R668 VSS.t23 VSS.n38 231.77
R669 VSS.t59 VSS.n8 231.77
R670 VSS.t49 VSS.n16 231.683
R671 VSS.t46 VSS.n148 231.683
R672 VSS.n152 VSS.t29 231.683
R673 VSS.n151 VSS.t26 231.683
R674 VSS.n105 VSS.t7 199.435
R675 VSS.n149 VSS.t3 199.435
R676 VSS.n207 VSS.t20 199.435
R677 VSS.n106 VSS.t13 194.475
R678 VSS.t5 VSS.n150 194.475
R679 VSS.n208 VSS.t18 194.475
R680 VSS.n148 VSS.n16 109.641
R681 VSS.n152 VSS.n151 71.44
R682 VSS.n106 VSS.n105 24.8059
R683 VSS.n150 VSS.n149 24.8059
R684 VSS.n208 VSS.n207 24.8059
R685 VSS.n93 VSS.n92 9.30555
R686 VSS.n166 VSS.t92 8.06917
R687 VSS.n166 VSS.t76 8.06917
R688 VSS.n163 VSS.t144 8.06917
R689 VSS.n163 VSS.t136 8.06917
R690 VSS.n162 VSS.t128 8.06917
R691 VSS.n162 VSS.t112 8.06917
R692 VSS.n156 VSS.t202 8.06917
R693 VSS.n156 VSS.t190 8.06917
R694 VSS.n155 VSS.t164 8.06917
R695 VSS.n155 VSS.t168 8.06917
R696 VSS.n219 VSS.t40 8.06917
R697 VSS.n219 VSS.t25 8.06917
R698 VSS.n166 VSS.t122 8.06917
R699 VSS.n166 VSS.t124 8.06917
R700 VSS.n163 VSS.t178 8.06917
R701 VSS.n163 VSS.t182 8.06917
R702 VSS.n162 VSS.t156 8.06917
R703 VSS.n162 VSS.t162 8.06917
R704 VSS.n156 VSS.t222 8.06917
R705 VSS.n156 VSS.t224 8.06917
R706 VSS.n155 VSS.t28 8.06917
R707 VSS.n155 VSS.t34 8.06917
R708 VSS.n219 VSS.t78 8.06917
R709 VSS.n219 VSS.t80 8.06917
R710 VSS.n81 VSS.t116 8.06917
R711 VSS.n80 VSS.t43 8.06917
R712 VSS.n87 VSS.t212 8.06917
R713 VSS.n79 VSS.t218 8.06917
R714 VSS.n201 VSS.t132 8.06917
R715 VSS.n175 VSS.t54 8.06917
R716 VSS.n9 VSS.t148 8.06917
R717 VSS.n171 VSS.t154 8.06917
R718 VSS.n198 VSS.t160 8.06917
R719 VSS.n198 VSS.t172 8.06917
R720 VSS.n196 VSS.t204 8.06917
R721 VSS.n196 VSS.t216 8.06917
R722 VSS.n195 VSS.t192 8.06917
R723 VSS.n195 VSS.t194 8.06917
R724 VSS.n191 VSS.t58 8.06917
R725 VSS.n191 VSS.t67 8.06917
R726 VSS.n190 VSS.t94 8.06917
R727 VSS.n190 VSS.t72 8.06917
R728 VSS.n188 VSS.t114 8.06917
R729 VSS.n188 VSS.t120 8.06917
R730 VSS.n99 VSS.t198 8.06917
R731 VSS.n69 VSS.t138 8.06917
R732 VSS.n39 VSS.t146 8.06917
R733 VSS.n65 VSS.t150 8.06917
R734 VSS.n62 VSS.t90 8.06917
R735 VSS.n62 VSS.t74 8.06917
R736 VSS.n60 VSS.t142 8.06917
R737 VSS.n60 VSS.t134 8.06917
R738 VSS.n59 VSS.t126 8.06917
R739 VSS.n59 VSS.t108 8.06917
R740 VSS.n55 VSS.t200 8.06917
R741 VSS.n55 VSS.t188 8.06917
R742 VSS.n54 VSS.t152 8.06917
R743 VSS.n54 VSS.t158 8.06917
R744 VSS.n52 VSS.t37 8.06917
R745 VSS.n52 VSS.t22 8.06917
R746 VSS.n132 VSS.t166 8.06917
R747 VSS.n110 VSS.t88 8.06917
R748 VSS.n47 VSS.t98 8.06917
R749 VSS.n46 VSS.t102 8.06917
R750 VSS.n26 VSS.t70 8.06917
R751 VSS.n25 VSS.t208 8.06917
R752 VSS.n32 VSS.t180 8.06917
R753 VSS.n24 VSS.t186 8.06917
R754 VSS.n76 VSS.t206 8.06917
R755 VSS.n76 VSS.t140 8.06917
R756 VSS.n73 VSS.t56 8.06917
R757 VSS.n73 VSS.t196 8.06917
R758 VSS.n72 VSS.t31 8.06917
R759 VSS.n72 VSS.t184 8.06917
R760 VSS.n143 VSS.t118 8.06917
R761 VSS.n143 VSS.t45 8.06917
R762 VSS.n142 VSS.t63 8.06917
R763 VSS.n142 VSS.t130 8.06917
R764 VSS.n139 VSS.t176 8.06917
R765 VSS.n139 VSS.t96 8.06917
R766 VSS.n76 VSS.t48 8.06917
R767 VSS.n76 VSS.t51 8.06917
R768 VSS.n73 VSS.t100 8.06917
R769 VSS.n73 VSS.t106 8.06917
R770 VSS.n72 VSS.t84 8.06917
R771 VSS.n72 VSS.t86 8.06917
R772 VSS.n143 VSS.t170 8.06917
R773 VSS.n143 VSS.t174 8.06917
R774 VSS.n142 VSS.t61 8.06917
R775 VSS.n142 VSS.t65 8.06917
R776 VSS.n139 VSS.t210 8.06917
R777 VSS.n139 VSS.t214 8.06917
R778 VSS.n182 VSS.t82 8.06917
R779 VSS.n183 VSS.t220 8.06917
R780 VSS.n212 VSS.t104 8.06917
R781 VSS.n5 VSS.t110 8.06917
R782 VSS.n119 VSS.n118 4.61205
R783 VSS.n126 VSS.n125 4.61205
R784 VSS.n116 VSS.n114 4.5005
R785 VSS.n123 VSS.n121 4.5005
R786 VSS.n112 VSS.n36 4.5005
R787 VSS.n112 VSS.n111 4.5005
R788 VSS.n130 VSS.n129 4.5005
R789 VSS.n131 VSS.n130 4.5005
R790 VSS.n113 VSS.t8 4.16278
R791 VSS.n120 VSS.t230 4.16278
R792 VSS.n118 VSS.n117 4.15984
R793 VSS.n125 VSS.n124 4.15984
R794 VSS.n127 VSS.n119 3.98482
R795 VSS.n113 VSS.t9 3.93054
R796 VSS.n120 VSS.t11 3.93054
R797 VSS.n116 VSS.n115 3.92774
R798 VSS.n123 VSS.n122 3.92774
R799 VSS.n88 VSS.t2 3.73318
R800 VSS.n91 VSS.n90 3.73318
R801 VSS.n88 VSS.t10 3.4916
R802 VSS.n91 VSS.n89 3.4916
R803 VSS.t117 VSS.n10 3.3605
R804 VSS.n84 VSS.t44 3.3605
R805 VSS.n86 VSS.t213 3.3605
R806 VSS.n96 VSS.t219 3.3605
R807 VSS.n200 VSS.t133 3.3605
R808 VSS.n204 VSS.t55 3.3605
R809 VSS.n174 VSS.t149 3.3605
R810 VSS.n170 VSS.t155 3.3605
R811 VSS.n98 VSS.t199 3.3605
R812 VSS.n102 VSS.t139 3.3605
R813 VSS.n68 VSS.t147 3.3605
R814 VSS.n64 VSS.t151 3.3605
R815 VSS.n135 VSS.t167 3.3605
R816 VSS.n109 VSS.t89 3.3605
R817 VSS.t99 VSS.n37 3.3605
R818 VSS.n50 VSS.t103 3.3605
R819 VSS.t71 VSS.n4 3.3605
R820 VSS.n29 VSS.t209 3.3605
R821 VSS.n31 VSS.t181 3.3605
R822 VSS.n35 VSS.t187 3.3605
R823 VSS.n186 VSS.t83 3.3605
R824 VSS.t221 VSS.n6 3.3605
R825 VSS.n211 VSS.t105 3.3605
R826 VSS.n215 VSS.t111 3.3605
R827 VSS.n127 VSS.n126 3.27473
R828 VSS.n114 VSS.n113 2.68012
R829 VSS.n121 VSS.n120 2.68012
R830 VSS.n34 VSS.n33 2.1005
R831 VSS.n28 VSS.n27 2.1005
R832 VSS.n49 VSS.n48 2.1005
R833 VSS.n134 VSS.n133 2.1005
R834 VSS.n67 VSS.n66 2.1005
R835 VSS.n101 VSS.n100 2.1005
R836 VSS.n214 VSS.n213 2.1005
R837 VSS.n185 VSS.n184 2.1005
R838 VSS.n173 VSS.n172 2.1005
R839 VSS.n203 VSS.n202 2.1005
R840 VSS.n95 VSS.n94 2.1005
R841 VSS.n83 VSS.n82 2.1005
R842 VSS.n128 VSS.n127 1.69669
R843 VSS.t44 VSS.n83 1.2605
R844 VSS.n83 VSS.t117 1.2605
R845 VSS.t219 VSS.n95 1.2605
R846 VSS.n95 VSS.t213 1.2605
R847 VSS.t55 VSS.n203 1.2605
R848 VSS.n203 VSS.t133 1.2605
R849 VSS.n173 VSS.t155 1.2605
R850 VSS.t149 VSS.n173 1.2605
R851 VSS.t139 VSS.n101 1.2605
R852 VSS.n101 VSS.t199 1.2605
R853 VSS.n67 VSS.t151 1.2605
R854 VSS.t147 VSS.n67 1.2605
R855 VSS.n134 VSS.t89 1.2605
R856 VSS.t167 VSS.n134 1.2605
R857 VSS.t103 VSS.n49 1.2605
R858 VSS.n49 VSS.t99 1.2605
R859 VSS.t209 VSS.n28 1.2605
R860 VSS.n28 VSS.t71 1.2605
R861 VSS.t187 VSS.n34 1.2605
R862 VSS.n34 VSS.t181 1.2605
R863 VSS.n185 VSS.t221 1.2605
R864 VSS.t83 VSS.n185 1.2605
R865 VSS.t111 VSS.n214 1.2605
R866 VSS.n214 VSS.t105 1.2605
R867 VSS.n11 VSS.t77 0.918039
R868 VSS.n12 VSS.t137 0.918039
R869 VSS.n13 VSS.t113 0.918039
R870 VSS.n154 VSS.t191 0.918039
R871 VSS.n0 VSS.t169 0.918039
R872 VSS.n3 VSS.t27 0.918039
R873 VSS.n167 VSS.t125 0.918039
R874 VSS.n164 VSS.t183 0.918039
R875 VSS.n160 VSS.t163 0.918039
R876 VSS.n157 VSS.t225 0.918039
R877 VSS.n1 VSS.t36 0.918039
R878 VSS.n217 VSS.t81 0.918039
R879 VSS.n176 VSS.t173 0.918039
R880 VSS.n177 VSS.t217 0.918039
R881 VSS.n178 VSS.t195 0.918039
R882 VSS.n179 VSS.t69 0.918039
R883 VSS.n180 VSS.t73 0.918039
R884 VSS.n181 VSS.t121 0.918039
R885 VSS.n40 VSS.t75 0.918039
R886 VSS.n41 VSS.t135 0.918039
R887 VSS.n42 VSS.t109 0.918039
R888 VSS.n43 VSS.t189 0.918039
R889 VSS.n44 VSS.t159 0.918039
R890 VSS.n45 VSS.t24 0.918039
R891 VSS.n70 VSS.t141 0.918039
R892 VSS.n71 VSS.t197 0.918039
R893 VSS.n17 VSS.t185 0.918039
R894 VSS.n21 VSS.t47 0.918039
R895 VSS.n22 VSS.t131 0.918039
R896 VSS.n23 VSS.t97 0.918039
R897 VSS.n77 VSS.t53 0.918039
R898 VSS.n74 VSS.t107 0.918039
R899 VSS.n18 VSS.t87 0.918039
R900 VSS.n144 VSS.t175 0.918039
R901 VSS.n140 VSS.t66 0.918039
R902 VSS.n137 VSS.t215 0.918039
R903 VSS.n11 VSS.t93 0.91749
R904 VSS.n12 VSS.t145 0.91749
R905 VSS.n13 VSS.t129 0.91749
R906 VSS.n154 VSS.t203 0.91749
R907 VSS.n0 VSS.t165 0.91749
R908 VSS.n3 VSS.t42 0.91749
R909 VSS.n167 VSS.t123 0.91749
R910 VSS.n164 VSS.t179 0.91749
R911 VSS.n160 VSS.t157 0.91749
R912 VSS.n157 VSS.t223 0.91749
R913 VSS.n1 VSS.t30 0.91749
R914 VSS.n217 VSS.t79 0.91749
R915 VSS.n176 VSS.t161 0.91749
R916 VSS.n177 VSS.t205 0.91749
R917 VSS.n178 VSS.t193 0.91749
R918 VSS.n179 VSS.t60 0.91749
R919 VSS.n180 VSS.t95 0.91749
R920 VSS.n181 VSS.t115 0.91749
R921 VSS.n40 VSS.t91 0.91749
R922 VSS.n41 VSS.t143 0.91749
R923 VSS.n42 VSS.t127 0.91749
R924 VSS.n43 VSS.t201 0.91749
R925 VSS.n44 VSS.t153 0.91749
R926 VSS.n45 VSS.t39 0.91749
R927 VSS.n70 VSS.t207 0.91749
R928 VSS.n71 VSS.t57 0.91749
R929 VSS.n17 VSS.t33 0.91749
R930 VSS.n21 VSS.t119 0.91749
R931 VSS.n22 VSS.t64 0.91749
R932 VSS.n23 VSS.t177 0.91749
R933 VSS.n77 VSS.t50 0.91749
R934 VSS.n74 VSS.t101 0.91749
R935 VSS.n18 VSS.t85 0.91749
R936 VSS.n144 VSS.t171 0.91749
R937 VSS.n140 VSS.t62 0.91749
R938 VSS.n137 VSS.t211 0.91749
R939 VSS.n138 VSS.n137 0.582999
R940 VSS.n141 VSS.n140 0.582999
R941 VSS.n145 VSS.n144 0.582999
R942 VSS.n19 VSS.n18 0.582999
R943 VSS.n75 VSS.n74 0.582999
R944 VSS.n78 VSS.n77 0.582999
R945 VSS.n138 VSS.n23 0.582999
R946 VSS.n141 VSS.n22 0.582999
R947 VSS.n145 VSS.n21 0.582999
R948 VSS.n19 VSS.n17 0.582999
R949 VSS.n75 VSS.n71 0.582999
R950 VSS.n78 VSS.n70 0.582999
R951 VSS.n51 VSS.n45 0.582999
R952 VSS.n53 VSS.n44 0.582999
R953 VSS.n56 VSS.n43 0.582999
R954 VSS.n58 VSS.n42 0.582999
R955 VSS.n61 VSS.n41 0.582999
R956 VSS.n63 VSS.n40 0.582999
R957 VSS.n187 VSS.n181 0.582999
R958 VSS.n189 VSS.n180 0.582999
R959 VSS.n192 VSS.n179 0.582999
R960 VSS.n194 VSS.n178 0.582999
R961 VSS.n197 VSS.n177 0.582999
R962 VSS.n199 VSS.n176 0.582999
R963 VSS.n218 VSS.n217 0.582999
R964 VSS.n2 VSS.n1 0.582999
R965 VSS.n158 VSS.n157 0.582999
R966 VSS.n161 VSS.n160 0.582999
R967 VSS.n165 VSS.n164 0.582999
R968 VSS.n168 VSS.n167 0.582999
R969 VSS.n218 VSS.n3 0.582999
R970 VSS.n2 VSS.n0 0.582999
R971 VSS.n158 VSS.n154 0.582999
R972 VSS.n161 VSS.n13 0.582999
R973 VSS.n165 VSS.n12 0.582999
R974 VSS.n168 VSS.n11 0.582999
R975 VSS.n92 VSS.n91 0.174974
R976 VSS.n119 VSS.n114 0.157683
R977 VSS.n126 VSS.n121 0.157683
R978 VSS.n92 VSS.n88 0.130788
R979 VSS.n104 VSS.n103 0.0886356
R980 VSS.n105 VSS.n104 0.0886356
R981 VSS.n57 VSS.n38 0.0886356
R982 VSS.n146 VSS.n20 0.0886356
R983 VSS.n20 VSS.n16 0.0886356
R984 VSS.n147 VSS.n146 0.0886356
R985 VSS.n148 VSS.n147 0.0886356
R986 VSS.n193 VSS.n8 0.0886356
R987 VSS.n206 VSS.n205 0.0886356
R988 VSS.n207 VSS.n206 0.0886356
R989 VSS.n85 VSS.n14 0.0886356
R990 VSS.n149 VSS.n14 0.0886356
R991 VSS.n159 VSS.n153 0.0886356
R992 VSS.n153 VSS.n152 0.0886356
R993 VSS.n159 VSS.n7 0.0886356
R994 VSS.n151 VSS.n7 0.0886356
R995 VSS.n108 VSS.n107 0.0871667
R996 VSS.n107 VSS.n106 0.0871667
R997 VSS.n30 VSS.n15 0.0871667
R998 VSS.n150 VSS.n15 0.0871667
R999 VSS.n210 VSS.n209 0.0871667
R1000 VSS.n209 VSS.n208 0.0871667
R1001 VSS.n198 VSS.n197 0.0390622
R1002 VSS.n189 VSS.n188 0.0390622
R1003 VSS.n62 VSS.n61 0.0385696
R1004 VSS.n53 VSS.n52 0.0385696
R1005 VSS.n196 VSS.n195 0.0371211
R1006 VSS.n191 VSS.n190 0.0371211
R1007 VSS.n60 VSS.n59 0.0366533
R1008 VSS.n55 VSS.n54 0.0366533
R1009 VSS.n65 VSS.n64 0.0341
R1010 VSS.n66 VSS.n65 0.0341
R1011 VSS.n66 VSS.n39 0.0341
R1012 VSS.n68 VSS.n39 0.0341
R1013 VSS.n102 VSS.n69 0.0341
R1014 VSS.n100 VSS.n69 0.0341
R1015 VSS.n100 VSS.n99 0.0341
R1016 VSS.n99 VSS.n98 0.0341
R1017 VSS.n171 VSS.n170 0.0341
R1018 VSS.n172 VSS.n171 0.0341
R1019 VSS.n172 VSS.n9 0.0341
R1020 VSS.n174 VSS.n9 0.0341
R1021 VSS.n204 VSS.n175 0.0341
R1022 VSS.n202 VSS.n175 0.0341
R1023 VSS.n202 VSS.n201 0.0341
R1024 VSS.n201 VSS.n200 0.0341
R1025 VSS.n96 VSS.n79 0.0341
R1026 VSS.n94 VSS.n79 0.0341
R1027 VSS.n87 VSS.n86 0.0341
R1028 VSS.n84 VSS.n80 0.0341
R1029 VSS.n82 VSS.n80 0.0341
R1030 VSS.n82 VSS.n81 0.0341
R1031 VSS.n81 VSS.n10 0.0341
R1032 VSS.n187 VSS.n186 0.0302339
R1033 VSS.n194 VSS.n193 0.0301981
R1034 VSS.n51 VSS.n50 0.0301505
R1035 VSS.n200 VSS.n199 0.0300328
R1036 VSS.n64 VSS.n63 0.0299989
R1037 VSS.n58 VSS.n57 0.0298187
R1038 VSS.n35 VSS.n24 0.0294988
R1039 VSS.n33 VSS.n24 0.0294988
R1040 VSS.n33 VSS.n32 0.0294988
R1041 VSS.n32 VSS.n31 0.0294988
R1042 VSS.n29 VSS.n25 0.0294988
R1043 VSS.n27 VSS.n25 0.0294988
R1044 VSS.n27 VSS.n26 0.0294988
R1045 VSS.n26 VSS.n4 0.0294988
R1046 VSS.n50 VSS.n46 0.0294988
R1047 VSS.n48 VSS.n46 0.0294988
R1048 VSS.n48 VSS.n47 0.0294988
R1049 VSS.n47 VSS.n37 0.0294988
R1050 VSS.n110 VSS.n109 0.0294988
R1051 VSS.n133 VSS.n110 0.0294988
R1052 VSS.n133 VSS.n132 0.0294988
R1053 VSS.n215 VSS.n5 0.0294988
R1054 VSS.n213 VSS.n5 0.0294988
R1055 VSS.n213 VSS.n212 0.0294988
R1056 VSS.n212 VSS.n211 0.0294988
R1057 VSS.n183 VSS.n6 0.0294988
R1058 VSS.n184 VSS.n183 0.0294988
R1059 VSS.n184 VSS.n182 0.0294988
R1060 VSS.n186 VSS.n182 0.0294988
R1061 VSS.n98 VSS.n97 0.02738
R1062 VSS.n170 VSS.n169 0.02738
R1063 VSS.n97 VSS.n96 0.02738
R1064 VSS.n169 VSS.n10 0.02738
R1065 VSS.n128 VSS.n112 0.0255051
R1066 VSS.n136 VSS.n35 0.0236991
R1067 VSS.n216 VSS.n4 0.0236991
R1068 VSS.n136 VSS.n135 0.0236991
R1069 VSS.n216 VSS.n215 0.0236991
R1070 VSS.n94 VSS.n93 0.022805
R1071 VSS.n130 VSS.n128 0.0215309
R1072 VSS.n193 VSS.n192 0.0203634
R1073 VSS.n57 VSS.n56 0.0201097
R1074 VSS.n103 VSS.n102 0.01994
R1075 VSS.n205 VSS.n204 0.01994
R1076 VSS.n85 VSS.n84 0.01994
R1077 VSS.n199 VSS.n198 0.0196517
R1078 VSS.n197 VSS.n196 0.0196517
R1079 VSS.n195 VSS.n194 0.0196517
R1080 VSS.n192 VSS.n191 0.0196517
R1081 VSS.n190 VSS.n189 0.0196517
R1082 VSS.n188 VSS.n187 0.0196517
R1083 VSS.n166 VSS.n165 0.0194273
R1084 VSS.n63 VSS.n62 0.019407
R1085 VSS.n61 VSS.n60 0.019407
R1086 VSS.n59 VSS.n58 0.019407
R1087 VSS.n56 VSS.n55 0.019407
R1088 VSS.n54 VSS.n53 0.019407
R1089 VSS.n52 VSS.n51 0.019407
R1090 VSS.n76 VSS.n75 0.0189267
R1091 VSS.n141 VSS.n139 0.0189267
R1092 VSS.n163 VSS.n162 0.0184746
R1093 VSS.n156 VSS.n155 0.0184746
R1094 VSS.n31 VSS.n30 0.0183136
R1095 VSS.n108 VSS.n37 0.0183136
R1096 VSS.n211 VSS.n210 0.0183136
R1097 VSS.n73 VSS.n72 0.0179991
R1098 VSS.n143 VSS.n142 0.0179991
R1099 VSS.n103 VSS.n68 0.01514
R1100 VSS.n205 VSS.n174 0.01514
R1101 VSS.n86 VSS.n85 0.01514
R1102 VSS.n161 VSS.n159 0.0150766
R1103 VSS.n146 VSS.n19 0.014691
R1104 VSS.n135 VSS.n36 0.0141709
R1105 VSS VSS.n2 0.0139016
R1106 VSS.n129 VSS.n111 0.0132388
R1107 VSS.n93 VSS.n87 0.0127708
R1108 VSS.n30 VSS.n29 0.0120995
R1109 VSS.n109 VSS.n108 0.0120995
R1110 VSS.n210 VSS.n6 0.0120995
R1111 VSS.n159 VSS.n158 0.0102495
R1112 VSS.n146 VSS.n145 0.00999158
R1113 VSS.n168 VSS.n166 0.00990014
R1114 VSS.n165 VSS.n163 0.00990014
R1115 VSS.n162 VSS.n161 0.00990014
R1116 VSS.n158 VSS.n156 0.00990014
R1117 VSS.n155 VSS.n2 0.00990014
R1118 VSS.n219 VSS.n218 0.00990014
R1119 VSS.n78 VSS.n76 0.00965149
R1120 VSS.n75 VSS.n73 0.00965149
R1121 VSS.n72 VSS.n19 0.00965149
R1122 VSS.n145 VSS.n143 0.00965149
R1123 VSS.n142 VSS.n141 0.00965149
R1124 VSS.n139 VSS.n138 0.00965149
R1125 VSS VSS.n219 0.00602576
R1126 VSS.n118 VSS.n116 0.00523684
R1127 VSS.n125 VSS.n123 0.00523684
R1128 VSS.n218 VSS.n216 0.00370748
R1129 VSS.n138 VSS.n136 0.00362264
R1130 VSS.n132 VSS.n131 0.00288205
R1131 VSS.n169 VSS.n168 0.00180205
R1132 VSS.n97 VSS.n78 0.00176761
R1133 VSS.n131 VSS.n111 0.000603567
R1134 VSS.n129 VSS.n36 0.000603567
R1135 a_n160_6615.t10 a_n160_6615.t3 12.7127
R1136 a_n160_6615.t10 a_n160_6615.t6 10.2828
R1137 a_n160_6615.t10 a_n160_6615.t0 10.2828
R1138 a_n160_6615.t10 a_n160_6615.t14 10.2828
R1139 a_n160_6615.t10 a_n160_6615.t15 10.2828
R1140 a_n160_6615.t10 a_n160_6615.t20 10.1333
R1141 a_n160_6615.t10 a_n160_6615.t24 10.1333
R1142 a_n160_6615.t10 a_n160_6615.t2 10.1333
R1143 a_n160_6615.t10 a_n160_6615.t4 10.1333
R1144 a_n160_6615.t10 a_n160_6615.t11 9.72545
R1145 a_n160_6615.t10 a_n160_6615.t17 9.57156
R1146 a_n160_6615.t10 a_n160_6615.t13 9.57156
R1147 a_n160_6615.t10 a_n160_6615.t19 9.57156
R1148 a_n160_6615.t10 a_n160_6615.t16 9.57156
R1149 a_n160_6615.t10 a_n160_6615.t23 9.57156
R1150 a_n160_6615.t10 a_n160_6615.t21 9.57156
R1151 a_n160_6615.t10 a_n160_6615.t25 9.57156
R1152 a_n160_6615.t10 a_n160_6615.t22 9.57156
R1153 a_n160_6615.t11 a_n160_6615.n0 8.02945
R1154 a_n160_6615.t10 a_n160_6615.n1 8.02708
R1155 a_n160_6615.t10 a_n160_6615.n2 7.90829
R1156 a_n160_6615.n3 a_n160_6615.t10 7.90829
R1157 a_n160_6615.t10 a_n160_6615.t5 7.41776
R1158 a_11579_648.n1 a_11579_648.t7 10.2515
R1159 a_11579_648.n1 a_11579_648.t3 10.2515
R1160 a_11579_648.n1 a_11579_648.t16 10.2515
R1161 a_11579_648.n1 a_11579_648.t13 10.2515
R1162 a_11579_648.n1 a_11579_648.t9 10.096
R1163 a_11579_648.n1 a_11579_648.t19 10.0935
R1164 a_11579_648.n1 a_11579_648.t5 10.0859
R1165 a_11579_648.n1 a_11579_648.t22 10.0808
R1166 a_11579_648.n1 a_11579_648.t23 9.53981
R1167 a_11579_648.n1 a_11579_648.t14 9.53981
R1168 a_11579_648.n1 a_11579_648.t24 9.53981
R1169 a_11579_648.n1 a_11579_648.t18 9.53981
R1170 a_11579_648.n1 a_11579_648.t15 9.53744
R1171 a_11579_648.n1 a_11579_648.t12 9.53744
R1172 a_11579_648.n1 a_11579_648.t21 9.53744
R1173 a_11579_648.n1 a_11579_648.t17 9.53744
R1174 a_11579_648.n1 a_11579_648.n0 8.41434
R1175 a_11579_648.n1 a_11579_648.n3 8.14082
R1176 a_11579_648.n0 a_11579_648.n4 8.13828
R1177 a_11579_648.t0 a_11579_648.n2 7.96115
R1178 a_11579_648.t0 a_11579_648.n5 7.94694
R1179 a_11579_648.t0 a_11579_648.n1 7.50666
R1180 a_11579_648.n0 a_11579_648.t10 7.48586
R1181 a_11579_648.n1 a_11579_648.t6 7.48333
R1182 a_12_588.t4 a_12_588.t2 21.6693
R1183 a_12_588.t3 a_12_588.t2 15.3476
R1184 ITN.n10 ITN.t2 6.53843
R1185 ITN.n2 ITN.t5 6.50376
R1186 ITN.n2 ITN.n1 5.97717
R1187 ITN.n8 ITN.n2 4.03666
R1188 ITN.n6 ITN.n4 3.89695
R1189 ITN.n3 ITN.t0 3.89695
R1190 ITN.n6 ITN.n5 3.73116
R1191 ITN.n3 ITN.t4 3.73116
R1192 ITN ITN.n0 3.653
R1193 ITN.n8 ITN.n7 3.39813
R1194 ITN.n10 ITN.n9 3.30288
R1195 ITN.n7 ITN.n3 2.58466
R1196 ITN ITN.n10 2.3283
R1197 ITN.n7 ITN.n6 2.22759
R1198 ITN.n9 ITN.n8 0.67025
R1199 ITN.n9 ITN 0.56225
R1200 a_5850_6555.n6 a_5850_6555.n1 10.2377
R1201 a_5850_6555.n5 a_5850_6555.n8 10.2108
R1202 a_5850_6555.n5 a_5850_6555.t5 9.99909
R1203 a_5850_6555.t0 a_5850_6555.n6 9.80443
R1204 a_5850_6555.n6 a_5850_6555.n10 9.55135
R1205 a_5850_6555.n0 a_5850_6555.t18 8.17385
R1206 a_5850_6555.n3 a_5850_6555.t22 8.17299
R1207 a_5850_6555.n3 a_5850_6555.t19 8.17134
R1208 a_5850_6555.n0 a_5850_6555.t16 8.16754
R1209 a_5850_6555.n1 a_5850_6555.t13 8.10567
R1210 a_5850_6555.n1 a_5850_6555.t15 8.10567
R1211 a_5850_6555.n3 a_5850_6555.t23 8.10567
R1212 a_5850_6555.n3 a_5850_6555.t21 8.10567
R1213 a_5850_6555.n1 a_5850_6555.t9 8.10567
R1214 a_5850_6555.n1 a_5850_6555.t12 8.10567
R1215 a_5850_6555.n0 a_5850_6555.t20 8.10567
R1216 a_5850_6555.n0 a_5850_6555.t17 8.10567
R1217 a_5850_6555.n7 a_5850_6555.t7 7.74799
R1218 a_5850_6555.n4 a_5850_6555.t3 7.73052
R1219 a_5850_6555.n7 a_5850_6555.n9 7.46478
R1220 a_5850_6555.n4 a_5850_6555.n11 7.1311
R1221 a_5850_6555.n5 a_5850_6555.n7 2.2505
R1222 a_5850_6555.n6 a_5850_6555.n4 2.2505
R1223 a_5850_6555.n1 a_5850_6555.t8 8.35731
R1224 a_5850_6555.n0 a_5850_6555.t10 8.38107
R1225 a_5850_6555.n1 a_5850_6555.t14 8.37583
R1226 a_5850_6555.n1 a_5850_6555.n0 4.35656
R1227 a_5850_6555.n6 a_5850_6555.n5 2.96863
R1228 a_5850_6555.n2 a_5850_6555.n1 1.0882
R1229 a_5850_6555.n2 a_5850_6555.n3 1.08408
R1230 a_5850_6555.n2 a_5850_6555.t11 8.66753
R1231 VA.n1 VA.t1 9.33982
R1232 VA VA.n1 7.46489
R1233 VA VA.n0 3.47265
R1234 VA.n1 VA 0.899326
R1235 a_5696_3730.t2 a_5696_3730.n0 10.3829
R1236 a_5696_3730.n0 a_5696_3730.t0 10.3566
R1237 a_5696_3730.n0 a_5696_3730.n2 10.0407
R1238 a_5696_3730.n0 a_5696_3730.n1 9.57605
R1239 a_5696_648.n0 a_5696_648.t0 10.6581
R1240 a_5696_648.t2 a_5696_648.n0 10.2346
R1241 a_5696_648.n0 a_5696_648.n2 9.5029
R1242 a_5696_648.n0 a_5696_648.n1 9.34796
R1243 VB.n1 VB.n0 9.24966
R1244 VB VB.n1 8.04195
R1245 VB VB.t1 3.46791
R1246 VB.n1 VB 1.01476
C0 ITN a_1816_3730# 0.04223f
C1 ITN IBN 1.68838f
C2 a_7622_1806# VDD 0.042519f
C3 IBN a_412_3730# 0.094151f
C4 VA IBP 0.271933f
C5 VDD a_12130_8547# 0.017204f
C6 VA a_7656_9713# 0.02829f
C7 a_1776_6615# VDD 0.05812f
C8 ITP VDD 2.69098f
C9 VDD a_370_7781# 0.062166f
C10 IBP a_13536_6615# 0.140064f
C11 IBP a_12130_7781# 0.093205f
C12 IBN a_1816_648# 0.146618f
C13 IBP a_13536_8547# 0.14146f
C14 VA VDD 1.47013f
C15 ITN a_412_1806# 0.056112f
C16 ITN a_1816_2572# 0.029143f
C17 ITP a_12130_8547# 0.039042f
C18 IBP VB 1.59009f
C19 VDD a_6250_9713# 0.021314f
C20 VDD a_13536_6615# 0.021515f
C21 VDD a_12130_7781# 0.017204f
C22 IBP a_6250_7781# 0.041194f
C23 VDD a_370_9713# 0.073724f
C24 IBN a_1816_3730# 0.063826f
C25 IBP a_7656_8547# 0.050814f
C26 a_370_8547# VDD 0.076387f
C27 IBP a_13536_7781# 0.060965f
C28 IBP a_7656_7781# 0.047571f
C29 VDD VB 1.72695f
C30 ITN a_412_648# 0.055873f
C31 a_7656_6615# VB 0.02829f
C32 ITN a_1816_1806# 0.042422f
C33 a_6218_1806# IBN 0.029151f
C34 ITP a_13536_6615# 0.042056f
C35 ITP a_12130_7781# 0.05261f
C36 a_12130_6615# VDD 0.029536f
C37 a_7622_2572# IBN 0.058572f
C38 IBP a_13536_9713# 0.05861f
C39 a_13536_7781# VDD 0.011958f
C40 ITP a_13536_8547# 0.029048f
C41 VDD a_6250_6615# 0.021515f
C42 IBP a_12130_9713# 0.09316f
C43 a_370_6615# VDD 0.073394f
C44 a_7622_648# IBN 0.041096f
C45 IBP a_6250_8547# 0.029183f
C46 IBP a_7656_9713# 0.021651f
C47 IBN a_412_1806# 0.094138f
C48 IBN a_1816_2572# 0.148015f
C49 ITN a_412_3730# 0.05592f
C50 IBN VDD 1.39949f
C51 VDD a_1776_7781# 0.046892f
C52 IBN a_6218_2572# 0.042325f
C53 VDD a_13536_9713# 0.024605f
C54 VDD a_12130_9713# 0.029536f
C55 VA VB 0.320841f
C56 IBP VDD 8.9594f
C57 a_12130_6615# ITP 0.05205f
C58 a_7656_9713# VDD 0.021314f
C59 a_13536_7781# ITP 0.042616f
C60 IBN a_7622_1806# 0.063642f
C61 a_6218_1806# VDD 0.042519f
C62 ITN a_1816_648# 0.042182f
C63 a_7622_2572# VDD 0.034176f
C64 VB a_6250_9713# 0.02829f
C65 VA a_6250_6615# 0.02829f
C66 VDD a_1776_9713# 0.05845f
C67 a_1776_8547# VDD 0.061113f
C68 IBN a_1816_1806# 0.065493f
C69 ITP a_13536_9713# 0.029004f
C70 ITP a_12130_9713# 0.038998f
C71 ITN a_412_2572# 0.042833f
C72 VDD a_6218_2572# 0.029136f
C73 IBP ITP 2.13747f
C74 a_7656_6615# VDD 0.021515f
.ends

