* Extracted by KLayout with GF180MCU LVS runset on : 05/04/2024 20:35

.SUBCKT Pass_tran VDD G D
M$1 D G VDD VDD pfet_03v3 L=1U W=16U AS=10.4P AD=6.72P PS=33.3U PD=16.84U
M$2 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$3 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$4 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$5 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$6 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$7 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$8 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$9 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$10 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$11 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$12 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$13 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$14 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$15 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$16 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$17 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$18 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$19 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$20 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$21 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$22 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$23 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$24 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$25 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$26 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$27 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$28 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$29 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$30 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$31 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$32 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$33 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$34 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$35 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$36 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$37 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$38 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$39 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$40 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$41 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$42 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$43 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$44 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$45 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$46 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$47 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$48 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$49 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$50 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=10.4P PS=16.84U PD=33.3U
M$51 D G VDD VDD pfet_03v3 L=1U W=16U AS=10.4P AD=6.72P PS=33.3U PD=16.84U
M$52 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$53 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$54 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$55 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$56 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$57 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$58 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$59 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$60 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$61 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$62 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$63 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$64 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$65 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$66 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$67 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$68 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$69 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$70 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$71 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$72 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$73 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$74 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$75 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$76 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$77 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$78 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$79 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$80 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$81 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$82 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$83 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$84 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$85 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$86 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$87 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$88 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$89 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$90 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$91 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$92 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$93 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$94 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$95 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$96 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$97 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$98 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$99 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$100 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=10.4P PS=16.84U PD=33.3U
M$101 D G VDD VDD pfet_03v3 L=1U W=16U AS=10.4P AD=6.72P PS=33.3U PD=16.84U
M$102 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$103 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$104 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$105 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$106 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$107 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$108 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$109 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$110 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$111 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$112 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$113 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$114 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$115 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$116 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$117 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$118 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$119 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$120 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$121 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$122 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$123 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$124 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$125 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$126 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$127 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$128 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$129 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$130 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$131 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$132 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$133 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$134 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$135 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$136 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$137 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$138 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$139 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$140 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$141 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$142 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$143 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$144 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$145 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$146 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$147 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$148 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$149 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$150 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=10.4P PS=16.84U PD=33.3U
M$151 D G VDD VDD pfet_03v3 L=1U W=16U AS=10.4P AD=6.72P PS=33.3U PD=16.84U
M$152 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$153 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$154 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$155 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$156 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$157 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$158 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$159 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$160 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$161 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$162 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$163 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$164 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$165 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$166 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$167 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$168 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$169 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$170 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$171 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$172 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$173 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$174 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$175 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$176 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$177 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$178 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$179 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$180 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$181 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$182 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$183 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$184 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$185 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$186 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$187 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$188 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$189 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$190 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$191 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$192 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$193 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$194 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$195 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$196 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$197 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$198 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$199 D G VDD VDD pfet_03v3 L=1U W=16U AS=6.72P AD=6.72P PS=16.84U PD=16.84U
M$200 VDD G D VDD pfet_03v3 L=1U W=16U AS=6.72P AD=10.4P PS=16.84U PD=33.3U
.ENDS Pass_tran
