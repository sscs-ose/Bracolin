* NGSPICE file created from Filter_TOP.ext - technology: gf180mcuD

.subckt Filter_TOP
X0 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3 a_118732_12343# PRbiased_net_5.IBP a_112452_9185# PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X7 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X8 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X9 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X10 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X11 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X12 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X13 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X14 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X15 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X16 a_29076_n27379# CM_n_net_0.IN a_28554_n28276# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X17 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X18 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X19 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X20 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X21 a_54966_3278# a_47184_10411# a_47356_3218# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X22 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X23 a_106972_n6007# a_106442_n7939# a_106442_n7939# PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X24 a_62154_n36281# CM_p_net_0.IN a_61624_n35376# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X25 a_47356_3218# a_47184_10411# a_53562_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X26 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X27 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X28 a_40734_n39838# CM_n_net_0.IN a_40174_n39838# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X29 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X30 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X31 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X32 a_118732_10411# PRbiased_net_5.IBP a_112452_9185# PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X33 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X34 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X35 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X36 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X37 a_112452_9185# PRbiased_net_5.IBP a_120138_11177# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X38 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X39 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X40 FC_top_0.AVDD FC_top_0.IREF a_n11312_n20927# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X41 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X42 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X43 PRbiased_net_0.VDD a_106442_n7939# a_106972_n6773# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X44 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X45 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X46 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X47 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X48 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X49 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X50 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X51 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X52 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X53 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X54 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X55 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X56 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X57 a_92469_4887# a_86091_10096# PRbiased_net_6.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X58 PRbiased_net_4.VDD a_27682_n7939# a_28212_n6007# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X59 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X60 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X61 a_34468_n39838# CM_n_net_0.IN a_33908_n39838# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X62 a_91947_6045# a_92101_8870# a_92501_12028# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X63 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X64 PRbiased_net_0.VDD a_106442_n7939# a_106972_n4841# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X65 FC_top_0.AVSS a_97830_n14221# a_98352_n14221# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X66 a_62154_n26431# CM_p_net_0.IN a_61624_n26431# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X67 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X68 a_57294_n26431# CM_p_net_0.IN a_56456_n26431# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X69 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X70 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X71 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X72 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X73 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X74 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X75 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X76 a_39421_3278# a_39421_3278# a_41347_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X77 a_43602_n22894# CM_n_net_0.IN a_43042_n21997# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X78 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X79 a_28212_n6773# a_27682_n7939# a_27682_n6773# PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X80 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X81 a_35902_n33559# CM_n_net_0.IN a_35342_n32662# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X82 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X83 a_n13565_n12405# a_n11312_n21934# a_5821_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X84 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X85 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X86 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X87 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X88 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X89 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X90 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X91 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X92 a_53040_n23716# CM_p_net_0.IN a_52732_n20096# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X93 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X94 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X95 a_68756_10862# a_66820_8930# PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X96 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X97 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X98 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X99 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X100 a_37336_n39838# CM_n_net_0.IN a_36776_n38941# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X101 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X102 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X103 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X104 a_28212_n4841# a_27682_n7939# a_27682_n6773# PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X105 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X106 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X107 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X108 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X109 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X110 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X111 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X112 FC_top_0.AVDD FC_top_0.IREF a_n11312_n21934# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X113 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X114 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X115 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X116 a_29636_n33559# CM_n_net_0.IN a_29076_n32662# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X117 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X118 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X119 a_97830_2963# a_86263_2903# a_99787_12028# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X120 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X121 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X122 a_52164_n25526# CM_p_net_0.IN a_51596_n25526# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X123 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X124 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X125 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X126 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X127 a_5821_n12405# a_n11312_n21934# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X128 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X129 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X130 a_5821_n12405# a_n11312_n21934# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X131 a_64128_n20096# CM_p_net_0.IN a_63560_n20096# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X132 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X133 a_58738_n23716# CM_p_net_0.IN a_58430_n20096# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X134 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X135 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X136 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X137 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X138 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X139 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X140 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X141 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X142 a_50758_n25526# CM_p_net_0.IN a_50228_n26431# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X143 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X144 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X145 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X146 a_114258_n6773# a_112452_n7999# FC_top_0.AVSS PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X147 a_99756_n13063# a_97830_n14221# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X148 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X149 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X150 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X151 a_29658_4436# a_27854_3218# PRbiased_net_9.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X152 a_92469_2963# a_86091_10096# a_91947_2963# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X153 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X154 a_33538_3278# a_33692_9185# a_34092_9245# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X155 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X156 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X157 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X158 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X159 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X160 a_114258_n4841# a_112452_n7999# a_112298_n13906# PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X161 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X162 FC_top_0.AVSS a_53194_9185# a_53594_11177# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X163 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X164 a_114224_4436# a_106442_10411# PRbiased_net_5.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X165 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X166 a_37336_n29173# CM_n_net_0.IN a_36776_n29173# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X167 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X168 a_49160_n13906# PRbiased_net_3.IBN PRbiased_net_3.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X169 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X170 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X171 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X172 PRbiased_net_4.IBP a_33692_n7999# a_35498_n6773# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X173 PRbiased_net_3.ITP PRbiased_net_3.IBP a_59474_n6773# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X174 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X175 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X176 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X177 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X178 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X179 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X180 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X181 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X182 a_62154_n34471# CM_p_net_0.IN a_61624_n34471# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X183 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X184 a_39972_9245# a_27854_3218# a_39421_3278# PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X185 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X186 a_57294_n34471# CM_p_net_0.IN a_56456_n34471# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X187 a_31070_n35353# CM_n_net_0.IN a_30510_n34456# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X188 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X189 a_57862_n27336# CM_p_net_0.IN a_57294_n27336# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X190 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X191 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X192 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X193 PRbiased_net_4.VA a_33692_n7999# a_35498_n4841# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X194 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X195 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X196 PRbiased_net_3.ITP PRbiased_net_3.IBP a_59474_n4841# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X197 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X198 a_106442_10411# a_106442_9245# a_108378_9245# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X199 a_47184_n6773# a_47184_n7939# a_49120_n7939# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X200 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X201 PRbiased_net_5.ITN a_106614_3218# a_107014_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X202 PRbiased_net_3.ITN a_47356_n13966# a_47756_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X203 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X204 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X205 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X206 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X207 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X208 a_56456_n27336# CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X209 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X210 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X211 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X212 a_31070_n24688# CM_n_net_0.IN a_30510_n23791# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X213 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X214 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X215 a_118703_n13906# a_118181_n13906# a_118181_n13906# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X216 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X217 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X218 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X219 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X220 a_33908_n28276# CM_n_net_0.IN a_33386_n29173# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X221 FC_top_0.AVDD FC_top_0.IREF a_n11312_n20927# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X222 a_54966_5202# a_47184_10411# PRbiased_net_8.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X223 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X224 a_52164_n33566# CM_p_net_0.IN a_51596_n33566# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X225 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X226 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X227 PRbiased_net_0.ITP a_106614_n13966# a_118732_n7939# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X228 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X229 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X230 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X231 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X232 a_53570_n21906# CM_p_net_0.IN a_52732_n21001# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X233 a_73230_8930# a_72830_8870# PRbiased_net_7.VA PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X234 a_29618_9245# a_27682_9245# PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X235 PRbiased_net_5.VA a_112452_9185# a_114258_12343# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X236 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X237 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X238 a_27682_9245# a_27854_3218# a_29658_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X239 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X240 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X241 a_n11312_n21934# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X242 a_40734_n38941# CM_n_net_0.IN a_40174_n38941# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X243 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X244 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X245 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X246 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X247 a_50758_n33566# CM_p_net_0.IN a_50228_n34471# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X248 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X249 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X250 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X251 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X252 PRbiased_net_5.IBP a_112452_9185# a_114258_10411# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X253 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X254 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X255 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X256 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X257 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X258 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X259 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X260 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X261 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X262 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X263 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X264 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X265 a_93873_n11139# a_86091_n7088# a_86263_n14281# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X266 a_64128_n21001# CM_p_net_0.IN a_63560_n21001# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X267 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X268 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X269 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X270 a_59268_n21906# CM_p_net_0.IN a_58430_n21001# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X271 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X272 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X273 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X274 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X275 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X276 a_34468_n38941# CM_n_net_0.IN a_33908_n38941# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X277 a_74602_n12297# a_66820_n7088# PRbiased_net_2.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X278 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X279 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X280 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X281 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X282 a_28254_6360# PRbiased_net_9.IBN a_27682_10411# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X283 a_118181_3278# a_118181_3278# a_120107_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X284 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X285 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X286 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X287 a_50758_n24621# CM_p_net_0.IN a_50228_n28241# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X288 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X289 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X290 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X291 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X292 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X293 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X294 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X295 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X296 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X297 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X298 a_37336_n24688# CM_n_net_0.IN a_36776_n24688# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X299 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X300 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X301 FC_top_0.AVDD FC_top_0.IREF a_n11312_n20927# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X302 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X303 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X304 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X305 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X306 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X307 PRbiased_net_2.IBN a_66820_n7088# a_73198_n13063# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X308 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X309 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X310 a_64966_n27336# CM_p_net_0.IN a_64128_n27336# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X311 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X312 a_40734_n29173# CM_n_net_0.IN a_40174_n29173# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X313 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X314 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X315 a_56456_n36281# CM_p_net_0.IN a_55926_n35376# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X316 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X317 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X318 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X319 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X320 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X321 a_27854_n13966# a_27682_n6773# a_34060_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X322 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X323 a_93907_n7088# a_92101_n8314# FC_top_0.AVSS PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X324 a_57862_n26431# CM_p_net_0.IN a_57294_n26431# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X325 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X326 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X327 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X328 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X329 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X330 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X331 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X332 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X333 a_55000_12343# a_53194_9185# a_53040_3278# PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X334 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X335 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X336 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X337 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X338 a_35342_n21997# CM_n_net_0.IN a_34468_n25585# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X339 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X340 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X341 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X342 a_34468_n29173# CM_n_net_0.IN a_33908_n29173# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X343 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X344 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X345 a_93907_n5156# a_92101_n8314# a_91947_n14221# PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X346 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X347 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X348 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X349 FC_top_0.AVDD FC_top_0.IREF a_n11312_n21934# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X350 PRbiased_net_1.VDD a_86091_n8254# a_86621_n7088# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X351 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X352 a_56456_n26431# CM_p_net_0.IN a_55926_n26431# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X353 FC_top_0.VOUT a_n11312_n21934# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X354 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X355 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X356 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X357 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X358 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X359 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X360 a_55000_10411# a_53194_9185# FC_top_0.AVSS PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X361 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X362 a_43042_n36250# CM_n_net_0.IN a_42168_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X363 FC_top_0.VOUT a_n11312_n21934# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X364 a_29618_12343# a_27682_9245# PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X365 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X366 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X367 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X368 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X369 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X370 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X371 PRbiased_net_8.VDD a_47184_9245# a_47714_12343# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X372 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X373 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X374 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X375 a_29076_n21997# CM_n_net_0.IN a_28202_n25585# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X376 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X377 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X378 a_n11312_n21934# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X379 PRbiased_net_1.VDD a_86091_n8254# a_86621_n5156# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X380 a_52164_n32661# CM_p_net_0.IN a_51596_n32661# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X381 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X382 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X383 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X384 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X385 a_52732_n25526# CM_p_net_0.IN a_52164_n25526# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X386 a_29618_10411# a_27682_9245# PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X387 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X388 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X389 PRbiased_net_8.VDD a_47184_9245# a_47714_10411# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X390 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X391 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X392 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X393 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X394 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X395 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X396 a_36776_n36250# CM_n_net_0.IN a_35902_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X397 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X398 a_43042_n25585# CM_n_net_0.IN a_42168_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X399 a_99787_n8254# PRbiased_net_1.IBP PRbiased_net_1.ITP PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X400 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X401 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X402 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X403 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X404 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X405 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X406 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X407 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X408 a_50758_n32661# CM_p_net_0.IN CM_p_net_0.OUT7 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X409 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X410 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X411 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X412 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X413 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X414 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X415 a_41608_n27379# CM_n_net_0.IN a_41086_n28276# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X416 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X417 PRbiased_net_1.IBN a_86091_n7088# a_92469_n13063# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X418 a_33908_n38044# CM_n_net_0.IN a_33386_n38044# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X419 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X420 a_35464_n12748# a_27682_n6773# PRbiased_net_4.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X421 a_n13565_n12405# a_n11312_n21934# a_5821_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X422 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X423 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X424 a_99787_n6322# PRbiased_net_1.IBP PRbiased_net_1.ITP PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X425 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X426 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X427 a_120138_n7939# PRbiased_net_0.IBP PRbiased_net_0.ITP PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X428 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X429 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X430 a_53040_6360# a_47184_10411# a_54966_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X431 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X432 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X433 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X434 a_64966_n36281# CM_p_net_0.IN a_64436_n35376# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X435 a_36776_n25585# CM_n_net_0.IN a_35902_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X436 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X437 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X438 a_40174_n36250# CM_n_net_0.IN CM_n_net_0.OUT12 FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X439 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X440 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X441 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X442 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X443 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X444 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X445 PRbiased_net_4.ITP PRbiased_net_4.IBP a_39972_n6773# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X446 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X447 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X448 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X449 a_57862_n34471# CM_p_net_0.IN a_57294_n34471# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X450 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X451 a_51596_n38996# CM_p_net_0.IN a_50758_n38996# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X452 a_58430_n27336# CM_p_net_0.IN a_57862_n27336# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X453 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X454 a_40734_n26482# CM_n_net_0.IN a_40174_n24688# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X455 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X456 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X457 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X458 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X459 a_73230_10096# a_72830_8870# PRbiased_net_7.IBP PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X460 a_106442_9245# a_106614_3218# a_108418_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X461 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X462 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X463 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X464 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X465 PRbiased_net_4.ITP PRbiased_net_4.IBP a_39972_n4841# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X466 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X467 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X468 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X469 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X470 a_40174_n25585# CM_n_net_0.IN CM_n_net_0.OUT6 FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X471 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X472 PRbiased_net_8.VB a_53194_9185# a_55000_9245# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X473 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X474 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X475 a_64966_n27336# CM_p_net_0.IN a_64128_n26431# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X476 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X477 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X478 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X479 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X480 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X481 a_53562_3278# a_47184_10411# a_53040_3278# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X482 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X483 a_118732_11177# a_106614_3218# a_118181_3278# PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X484 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X485 a_56456_n34471# CM_p_net_0.IN a_55926_n34471# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X486 a_47184_n6773# a_47184_n7939# a_49120_n6007# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X487 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X488 a_53040_n10824# a_47184_n6773# a_54966_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X489 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X490 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X491 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X492 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X493 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X494 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X495 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X496 a_34468_n26482# CM_n_net_0.IN a_33908_n24688# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X497 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X498 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X499 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X500 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X501 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X502 a_59445_n12748# a_58923_n13906# a_53194_n7999# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X503 a_74602_n14221# a_66820_n7088# a_66992_n14281# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X504 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X505 a_37336_n35353# CM_n_net_0.IN a_36776_n34456# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X506 FC_top_0.AVSS a_78559_n14221# a_79081_n13063# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X507 a_52732_n33566# CM_p_net_0.IN a_52164_n33566# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X508 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X509 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X510 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X511 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X512 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X513 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X514 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X515 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X516 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X517 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X518 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X519 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X520 a_108418_6360# a_106614_3218# PRbiased_net_5.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X521 a_35464_n10824# a_27682_n6773# a_27854_n13966# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X522 a_41347_n11982# a_39421_n13906# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X523 PRbiased_net_0.ITP a_106614_n13966# a_118732_n6007# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X524 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X525 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X526 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X527 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X528 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X529 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X530 FC_top_0.AVSS a_39421_3278# a_39943_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X531 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X532 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X533 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X534 a_37336_n24688# CM_n_net_0.IN a_36776_n23791# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X535 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X536 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X537 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X538 a_86091_n7088# PRbiased_net_1.IBN a_88067_n12297# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X539 a_39943_n13906# a_39421_n13906# a_39421_n13906# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X540 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X541 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X542 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X543 a_88027_n8254# a_86091_n8254# PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X544 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X545 PRbiased_net_6.VDD a_86091_8930# a_86621_8930# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X546 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X547 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X548 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X549 a_86091_10096# a_86091_8930# a_88027_8930# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X550 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X551 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X552 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X553 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X554 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X555 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X556 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X557 a_35902_n39838# CM_n_net_0.IN a_35342_n39838# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X558 a_33908_n33559# CM_n_net_0.IN a_33386_n33559# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X559 a_78559_2963# a_66992_2903# a_80516_10096# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X560 a_88027_n6322# a_86091_n8254# PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X561 PRbiased_net_5.IBN a_106442_10411# a_112820_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X562 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X563 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X564 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X565 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X566 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X567 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X568 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X569 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X570 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X571 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X572 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X573 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X574 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X575 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X576 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X577 PRbiased_net_7.ITP PRbiased_net_7.IBP a_79110_10096# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X578 a_64966_n37186# CM_p_net_0.IN a_64128_n34471# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X579 a_29636_n39838# CM_n_net_0.IN a_29076_n39838# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X580 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X581 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X582 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X583 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X584 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X585 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X586 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X587 a_59445_n10824# a_58923_n13906# a_53194_n7999# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X588 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X589 a_33908_n22894# CM_n_net_0.IN a_33386_n22894# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X590 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X591 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X592 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X593 a_92101_n8314# a_97830_n14221# a_99756_n12297# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X594 a_62992_n25526# CM_p_net_0.IN a_62154_n25526# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X595 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X596 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X597 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X598 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X599 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X600 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X601 a_43042_n35353# CM_n_net_0.IN a_42520_n37147# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X602 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X603 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X604 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X605 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X606 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X607 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X608 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X609 a_51596_n39901# CM_p_net_0.IN a_50758_n39901# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X610 FC_top_0.AVSS a_97830_n14221# a_98352_n13063# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X611 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X612 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X613 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X614 a_58430_n26431# CM_p_net_0.IN a_57862_n26431# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X615 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X616 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X617 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X618 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X619 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X620 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X621 a_112820_4436# a_106442_10411# PRbiased_net_5.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X622 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X623 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X624 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X625 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X626 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X627 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X628 a_36776_n35353# CM_n_net_0.IN a_36254_n37147# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X629 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X630 FC_top_0.AVDD FC_top_0.IREF a_n11312_n20927# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X631 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X632 a_5821_n12405# a_n11312_n21934# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X633 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X634 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X635 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X636 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X637 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X638 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X639 a_30510_n27379# CM_n_net_0.IN a_29988_n28276# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X640 PRbiased_net_8.VDD a_47184_10411# a_54966_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X641 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X642 a_n11312_n20927# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X643 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X644 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X645 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X646 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X647 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X648 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X649 a_73198_n11139# a_66820_n7088# a_72676_n11139# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X650 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X651 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X652 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X653 a_79110_n8254# a_66992_n14281# a_78559_n14221# PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X654 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X655 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X656 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X657 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X658 a_40734_n34456# CM_n_net_0.IN a_40174_n34456# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X659 a_52732_n32661# CM_p_net_0.IN a_52164_n32661# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X660 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X661 a_n11312_n21934# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X662 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X663 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X664 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X665 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X666 a_40174_n35353# CM_n_net_0.IN a_39652_n35353# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X667 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X668 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X669 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X670 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X671 FC_top_0.VOUT a_n11312_n21934# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X672 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X673 a_79110_n6322# a_66992_n14281# a_78559_n14221# PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X674 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X675 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X676 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X677 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X678 a_93873_6045# a_86091_10096# a_86263_2903# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X679 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X680 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X681 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X682 a_53562_5202# a_47184_10411# PRbiased_net_8.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X683 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X684 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X685 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X686 a_34468_n34456# CM_n_net_0.IN a_33908_n34456# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X687 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X688 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X689 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X690 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X691 a_40734_n23791# CM_n_net_0.IN a_40174_n23791# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X692 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X693 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X694 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X695 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X696 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X697 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X698 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X699 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X700 a_29658_3278# PRbiased_net_9.IBN PRbiased_net_9.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X701 PRbiased_net_9.ITN PRbiased_net_9.IBN a_28254_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X702 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X703 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X704 a_53570_n38996# CM_p_net_0.IN a_52732_n38996# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X705 a_27642_n27379# CM_n_net_0.IN a_27120_n27379# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X706 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X707 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X708 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X709 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X710 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X711 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X712 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X713 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X714 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X715 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X716 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X717 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X718 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X719 a_39943_6360# a_39421_3278# a_33692_9185# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X720 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X721 a_120138_n6007# PRbiased_net_0.IBP PRbiased_net_0.ITP PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X722 a_62992_n33566# CM_p_net_0.IN a_62154_n33566# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X723 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X724 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X725 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X726 a_93907_12028# a_92101_8870# a_91947_2963# PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X727 a_114224_3278# a_106442_10411# a_106614_3218# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X728 a_n11312_n20927# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X729 PRbiased_net_5.IBP a_112452_9185# a_114258_11177# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X730 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X731 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X732 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X733 a_49160_n12748# a_47356_n13966# PRbiased_net_3.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X734 a_34468_n23791# CM_n_net_0.IN a_33908_n23791# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X735 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X736 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X737 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X738 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X739 PRbiased_net_7.VDD a_66820_8930# a_67350_10096# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X740 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X741 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X742 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X743 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X744 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X745 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X746 a_58430_n34471# CM_p_net_0.IN a_57862_n34471# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X747 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X748 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X749 a_64128_n38996# CM_p_net_0.IN a_63560_n38996# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X750 PRbiased_net_6.VDD a_86091_8930# a_86621_12028# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X751 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X752 a_59268_n38996# CM_p_net_0.IN a_58430_n38996# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X753 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X754 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X755 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X756 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X757 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X758 a_86091_n7088# PRbiased_net_1.IBN a_88067_n14221# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X759 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X760 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X761 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X762 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X763 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X764 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X765 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X766 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X767 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X768 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X769 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X770 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X771 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X772 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X773 a_28202_n36250# CM_n_net_0.IN a_27642_n36250# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X774 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X775 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X776 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X777 a_118703_n12748# a_118181_n13906# a_112452_n7999# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X778 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X779 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X780 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X781 a_93873_4121# a_86091_10096# PRbiased_net_6.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X782 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X783 a_n13565_n11419# a_n11312_n21934# FC_top_0.VOUT FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X784 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X785 a_n13565_n11419# a_n11312_n21934# FC_top_0.VOUT FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X786 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X787 a_41608_n21997# CM_n_net_0.IN a_40734_n25585# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X788 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X789 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X790 a_35902_n39838# CM_n_net_0.IN a_35342_n38941# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X791 a_33908_n32662# CM_n_net_0.IN a_33386_n33559# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X792 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X793 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X794 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X795 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X796 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X797 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X798 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X799 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X800 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X801 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X802 a_28202_n25585# CM_n_net_0.IN a_27642_n25585# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X803 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X804 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X805 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X806 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X807 a_92101_n8314# a_97830_n14221# a_99756_n14221# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X808 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X809 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X810 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X811 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X812 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X813 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X814 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X815 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X816 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X817 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X818 a_49160_n10824# a_47356_n13966# PRbiased_net_3.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X819 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X820 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X821 a_92501_n8254# a_92101_n8314# PRbiased_net_1.VA PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X822 a_29636_n39838# CM_n_net_0.IN a_29076_n38941# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X823 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X824 a_55000_11177# a_53194_9185# FC_top_0.AVSS PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X825 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X826 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X827 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X828 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X829 a_108378_n6773# a_106442_n7939# PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X830 a_34092_n7939# a_33692_n7999# PRbiased_net_4.VA PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X831 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X832 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X833 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X834 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X835 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X836 a_30510_n37147# CM_n_net_0.IN a_29988_n37147# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X837 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X838 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X839 a_79081_n11139# a_78559_n14221# a_72830_n8314# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X840 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X841 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X842 a_92501_n6322# a_92101_n8314# PRbiased_net_1.IBP PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X843 a_53594_12343# a_53194_9185# PRbiased_net_8.VB PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X844 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X845 FC_top_0.AVDD FC_top_0.IREF a_n11312_n21934# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X846 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X847 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X848 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X849 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X850 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X851 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X852 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X853 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X854 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X855 a_29618_11177# a_27682_9245# PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X856 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X857 a_86621_8930# a_86091_8930# a_86091_8930# PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X858 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X859 a_108378_n4841# a_106442_n7939# PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X860 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X861 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X862 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X863 PRbiased_net_8.VDD a_47184_9245# a_47714_11177# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X864 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X865 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X866 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X867 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X868 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X869 CM_p_net_0.VDD CM_p_net_0.IN a_52732_n39901# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X870 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X871 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X872 a_35902_n29173# CM_n_net_0.IN a_35342_n29173# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X873 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X874 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X875 a_27682_n7939# a_27682_n7939# a_29618_n6773# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X876 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X877 a_53594_10411# a_53194_9185# PRbiased_net_8.IBP PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X878 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X879 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X880 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X881 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X882 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X883 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X884 a_30510_n26482# CM_n_net_0.IN a_29988_n26482# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X885 a_118703_n10824# a_118181_n13906# a_112452_n7999# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X886 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X887 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X888 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X889 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X890 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X891 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X892 a_62992_n32661# CM_p_net_0.IN a_62154_n32661# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X893 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X894 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X895 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X896 a_63560_n25526# CM_p_net_0.IN a_62992_n25526# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X897 PRbiased_net_8.VDD a_47184_9245# a_47714_9245# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X898 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X899 a_51596_n38091# CM_p_net_0.IN a_50758_n38091# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X900 FC_top_0.AVSS a_n11312_n20927# a_n11312_n20927# FC_top_0.AVSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X901 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X902 a_27682_n7939# a_27682_n7939# a_29618_n4841# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X903 a_58923_n13906# a_47356_n13966# a_60880_n6773# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X904 a_99787_n7088# a_86263_n14281# PRbiased_net_1.ITP PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X905 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X906 PRbiased_net_4.IBN a_27682_n6773# a_34060_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X907 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X908 a_86663_n11139# PRbiased_net_1.IBN a_86091_n7088# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X909 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X910 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X911 a_64128_n39901# CM_p_net_0.IN a_63560_n39901# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X912 a_29636_n29173# CM_n_net_0.IN a_29076_n29173# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X913 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X914 PRbiased_net_2.VB a_72830_n8314# a_74636_n8254# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X915 CM_p_net_0.VDD CM_p_net_0.IN a_58430_n39901# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X916 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X917 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X918 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X919 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X920 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X921 a_58923_n13906# a_47356_n13966# a_60880_n4841# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X922 a_27642_n37147# CM_n_net_0.IN a_27120_n38044# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X923 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X924 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X925 a_99787_n5156# a_86263_n14281# PRbiased_net_1.ITP PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X926 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X927 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X928 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X929 a_n11312_n20927# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X930 a_72830_8870# PRbiased_net_7.IBP a_80516_8930# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X931 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X932 a_29658_5202# PRbiased_net_9.IBN PRbiased_net_9.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X933 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X934 PRbiased_net_2.IBP a_72830_n8314# a_74636_n6322# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X935 a_108418_n13906# PRbiased_net_0.IBN PRbiased_net_0.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X936 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X937 PRbiased_net_8.ITN PRbiased_net_8.IBN a_47756_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X938 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X939 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X940 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X941 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X942 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X943 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X944 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X945 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X946 PRbiased_net_5.ITN PRbiased_net_5.IBN a_107014_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X947 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X948 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X949 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X950 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X951 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X952 a_114224_5202# a_106442_10411# PRbiased_net_5.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X953 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X954 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X955 a_106442_9245# a_106442_9245# a_108378_12343# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X956 a_27642_n26482# CM_n_net_0.IN a_27120_n27379# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X957 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X958 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X959 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X960 a_112452_n7999# PRbiased_net_0.IBP a_120138_n7939# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X961 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X962 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X963 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X964 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X965 a_98352_n11139# a_97830_n14221# a_92101_n8314# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X966 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X967 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X968 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X969 a_54966_6360# a_47184_10411# a_47356_3218# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X970 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X971 a_106442_9245# a_106442_9245# a_108378_10411# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X972 a_51596_n31756# CM_p_net_0.IN a_50758_n31756# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X973 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X974 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X975 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X976 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X977 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X978 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X979 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X980 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X981 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X982 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X983 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X984 a_73230_10862# a_72830_8870# PRbiased_net_7.IBP PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X985 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X986 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X987 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X988 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X989 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X990 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X991 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X992 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X993 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X994 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X995 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X996 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X997 a_93873_4887# a_86091_10096# PRbiased_net_6.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X998 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X999 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1000 a_120107_n13906# a_118181_n13906# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1001 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1002 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1003 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1004 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1005 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1006 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1007 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1008 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1009 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1010 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1011 a_27854_n13966# a_27682_n6773# a_34060_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1012 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1013 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1014 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1015 a_51596_n22811# CM_p_net_0.IN a_50758_n22811# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1016 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1017 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1018 a_93873_n12297# a_86091_n7088# PRbiased_net_1.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1019 a_63560_n33566# CM_p_net_0.IN a_62992_n33566# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1020 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1021 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1022 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1023 a_28202_n37147# CM_n_net_0.IN a_27642_n35353# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1024 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1025 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1026 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1027 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1028 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1029 a_30510_n21997# CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1030 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1031 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1032 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1033 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1034 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1035 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1036 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1037 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1038 a_88027_n7088# a_86091_n8254# PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1039 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1040 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1041 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1042 a_n11312_n21934# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1043 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1044 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1045 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1046 a_49120_12343# a_47184_9245# PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1047 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1048 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1049 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1050 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1051 PRbiased_net_3.VDD a_47184_n6773# a_54966_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1052 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1053 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1054 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1055 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1056 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1057 a_88027_n5156# a_86091_n8254# PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1058 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1059 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1060 a_74602_n13063# a_66820_n7088# PRbiased_net_2.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1061 a_43602_n29173# CM_n_net_0.IN a_43042_n28276# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1062 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1063 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1064 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1065 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1066 a_49120_10411# a_47184_9245# PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1067 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1068 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1069 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1070 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1071 a_72830_8870# PRbiased_net_7.IBP a_80516_10862# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1072 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1073 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1074 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1075 a_93873_2963# a_86091_10096# a_86263_2903# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1076 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1077 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1078 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1079 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1080 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1081 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1082 a_53040_n13906# a_53194_n7999# a_53594_n7939# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1083 a_27642_n21997# CM_n_net_0.IN a_27120_n22894# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1084 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1085 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1086 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1087 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1088 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1089 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1090 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1091 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1092 a_53570_n24621# CM_p_net_0.IN a_53040_n23716# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1093 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1094 PRbiased_net_7.ITP a_66992_2903# a_79110_10862# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1095 a_33538_n10824# a_27682_n6773# a_35464_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1096 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1097 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1098 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1099 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1100 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1101 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1102 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1103 FC_top_0.AVSS a_n11312_n20927# a_n11312_n20927# FC_top_0.AVSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X1104 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1105 a_91947_2963# a_86091_10096# a_93873_6045# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1106 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1107 a_39943_n12748# a_39421_n13906# a_33692_n7999# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1108 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1109 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1110 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1111 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1112 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1113 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1114 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1115 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1116 a_112852_n6773# a_112452_n7999# PRbiased_net_0.IBP PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1117 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1118 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1119 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1120 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1121 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1122 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1123 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1124 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1125 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1126 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1127 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1128 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1129 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1130 PRbiased_net_9.ITP a_27854_3218# a_39972_9245# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1131 a_34092_n6007# a_33692_n7999# PRbiased_net_4.IBP PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1132 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1133 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1134 a_106614_3218# a_106442_10411# a_112820_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1135 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1136 a_59268_n24621# CM_p_net_0.IN a_58738_n23716# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1137 FC_top_0.AVDD FC_top_0.IREF a_n11312_n21934# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1138 a_112852_n4841# a_112452_n7999# PRbiased_net_0.VB PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1139 a_53570_n38996# CM_p_net_0.IN a_52732_n38091# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1140 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1141 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1142 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1143 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1144 a_79110_n7088# PRbiased_net_2.IBP a_72830_n8314# PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1145 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1146 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1147 FC_top_0.AVSS a_33692_n7999# a_34092_n6773# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1148 a_53040_n13906# a_47184_n6773# a_54966_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1149 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1150 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1151 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1152 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1153 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1154 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1155 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1156 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1157 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1158 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1159 a_63560_n32661# CM_p_net_0.IN a_62992_n32661# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1160 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1161 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1162 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1163 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1164 a_67350_10096# a_66820_8930# a_66820_10096# PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1165 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1166 a_79110_n5156# PRbiased_net_2.IBP a_72830_n8314# PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1167 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1168 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1169 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1170 a_33538_n10824# a_33692_n7999# a_34092_n4841# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1171 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1172 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1173 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1174 FC_top_0.AVSS a_58923_n13906# a_59445_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1175 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X1176 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1177 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1178 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1179 a_64128_n38091# CM_p_net_0.IN a_63560_n38091# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1180 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1181 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1182 a_59268_n38996# CM_p_net_0.IN a_58430_n38091# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1183 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1184 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1185 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1186 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1187 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1188 PRbiased_net_5.VB a_112452_9185# a_114258_9245# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1189 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1190 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1191 a_112820_3278# a_106442_10411# a_112298_3278# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1192 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1193 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1194 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1195 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1196 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1197 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1198 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1199 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1200 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1201 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1202 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1203 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1204 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1205 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1206 PRbiased_net_6.VDD a_86091_10096# a_93873_4121# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1207 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1208 a_39943_n10824# a_39421_n13906# a_33692_n7999# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1209 a_35902_n34456# CM_n_net_0.IN a_35342_n34456# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1210 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1211 a_120138_9245# PRbiased_net_5.IBP PRbiased_net_5.ITP PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1212 a_93873_n14221# a_86091_n7088# a_86263_n14281# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1213 a_53040_n35376# CM_p_net_0.IN a_52732_n31756# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1214 a_112298_6360# a_112452_9185# a_112852_12343# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1215 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1216 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1217 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1218 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1219 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1220 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1221 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1222 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1223 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1224 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1225 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1226 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1227 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1228 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1229 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1230 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1231 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1232 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1233 a_29636_n34456# CM_n_net_0.IN a_29076_n34456# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1234 PRbiased_net_7.VDD a_66820_8930# a_67350_10862# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1235 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1236 FC_top_0.AVSS a_112452_9185# a_112852_10411# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1237 a_112452_n7999# PRbiased_net_0.IBP a_120138_n6007# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1238 a_35902_n23791# CM_n_net_0.IN a_35342_n23791# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1239 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1240 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1241 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1242 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1243 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1244 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1245 a_29658_n13906# PRbiased_net_4.IBN PRbiased_net_4.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1246 a_64128_n31756# CM_p_net_0.IN a_63560_n31756# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1247 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1248 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1249 a_41378_n6773# a_27854_n13966# PRbiased_net_4.ITP PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1250 a_35464_n11982# a_27682_n6773# PRbiased_net_4.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1251 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1252 a_53570_n25526# CM_p_net_0.IN a_52732_n22811# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1253 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1254 a_58738_n35376# CM_p_net_0.IN a_58430_n31756# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1255 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1256 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1257 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1258 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1259 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1260 a_43602_n38044# CM_n_net_0.IN a_43042_n38044# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1261 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1262 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1263 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1264 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1265 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1266 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1267 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1268 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1269 a_29636_n23791# CM_n_net_0.IN a_29076_n23791# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1270 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1271 a_41378_n4841# a_27854_n13966# PRbiased_net_4.ITP PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1272 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1273 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1274 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1275 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1276 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1277 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1278 a_99787_12028# a_86263_2903# PRbiased_net_6.ITP PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1279 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1280 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1281 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1282 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1283 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1284 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1285 a_33908_n39838# CM_n_net_0.IN a_33386_n39838# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1286 a_64128_n22811# CM_p_net_0.IN a_63560_n22811# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1287 a_60880_9245# PRbiased_net_8.IBP PRbiased_net_8.ITP PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1288 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1289 a_59268_n25526# CM_p_net_0.IN a_58430_n22811# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1290 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1291 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1292 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1293 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1294 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1295 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1296 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1297 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1298 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1299 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1300 a_92101_8870# PRbiased_net_6.IBP a_99787_8930# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1301 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1302 a_62154_n37186# CM_p_net_0.IN a_61624_n38091# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1303 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1304 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1305 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1306 a_57294_n37186# CM_p_net_0.IN a_56456_n37186# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1307 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1308 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1309 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1310 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1311 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1312 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1313 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1314 a_92501_n7088# a_92101_n8314# PRbiased_net_1.IBP PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1315 a_29636_n38044# CM_n_net_0.IN a_30510_n36250# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1316 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1317 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1318 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1319 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1320 a_86091_n8254# a_86263_n14281# a_88067_n13063# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1321 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1322 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1323 a_60880_n6773# a_47356_n13966# PRbiased_net_3.ITP PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1324 a_n11312_n21934# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1325 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1326 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1327 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1328 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1329 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1330 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1331 a_27682_10411# a_27682_9245# a_29618_9245# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1332 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1333 a_59445_n11982# a_58923_n13906# a_58923_n13906# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1334 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1335 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1336 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1337 a_92501_n5156# a_92101_n8314# PRbiased_net_1.VB PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1338 a_53594_11177# a_53194_9185# PRbiased_net_8.IBP PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1339 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1340 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1341 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1342 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1343 a_62154_n28241# CM_p_net_0.IN a_61624_n28241# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1344 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1345 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1346 a_60880_n4841# a_47356_n13966# PRbiased_net_3.ITP PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1347 a_35342_n28276# CM_n_net_0.IN a_34820_n28276# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1348 a_35498_n6773# a_33692_n7999# FC_top_0.AVSS PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1349 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1350 a_57294_n28241# CM_p_net_0.IN a_56456_n28241# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1351 PRbiased_net_5.IBN a_106442_10411# a_112820_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1352 a_59474_n6773# PRbiased_net_3.IBP a_53194_n7999# PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1353 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1354 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1355 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1356 a_29636_n27379# CM_n_net_0.IN a_30510_n25585# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1357 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1358 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1359 FC_top_0.AVSS a_58923_3278# a_59445_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1360 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1361 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1362 a_39421_3278# a_27854_3218# a_41378_12343# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1363 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1364 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1365 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1366 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1367 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1368 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1369 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1370 FC_top_0.AVDD FC_top_0.IREF a_n11312_n20927# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1371 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1372 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1373 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1374 FC_top_0.AVSS a_92101_8870# a_92501_10096# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1375 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1376 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1377 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1378 a_35498_n4841# a_33692_n7999# a_33538_n13906# PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1379 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1380 a_59474_n4841# PRbiased_net_3.IBP a_53194_n7999# PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1381 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1382 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1383 FC_top_0.AVSS a_53194_n7999# a_53594_n6007# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1384 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1385 a_53040_3278# a_47184_10411# a_54966_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1386 a_80516_n8254# PRbiased_net_2.IBP PRbiased_net_2.ITP PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1387 a_97830_n14221# a_97830_n14221# a_99756_n13063# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1388 a_29076_n28276# CM_n_net_0.IN a_28554_n28276# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1389 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1390 a_112298_n10824# a_106442_n6773# a_114224_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1391 a_39421_3278# a_27854_3218# a_41378_10411# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1392 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1393 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1394 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1395 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1396 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1397 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1398 PRbiased_net_2.IBP a_72830_n8314# a_74636_n7088# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1399 a_73198_n12297# a_66820_n7088# PRbiased_net_2.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1400 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1401 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1402 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1403 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1404 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1405 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1406 a_52164_n27336# CM_p_net_0.IN a_51596_n27336# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1407 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1408 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1409 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1410 a_72676_n14221# a_66820_n7088# a_74602_n11139# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1411 PRbiased_net_6.VDD a_86091_10096# a_93873_4887# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1412 a_112820_5202# a_106442_10411# PRbiased_net_5.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1413 a_80516_n6322# PRbiased_net_2.IBP PRbiased_net_2.ITP PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1414 a_43602_n33559# CM_n_net_0.IN a_43042_n33559# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1415 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1416 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1417 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1418 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1419 a_72676_n14221# a_72830_n8314# a_73230_n8254# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1420 PRbiased_net_2.VA a_72830_n8314# a_74636_n5156# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1421 a_118732_n7939# a_106614_n13966# a_118181_n13906# PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1422 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1423 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1424 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1425 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1426 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1427 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1428 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1429 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1430 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1431 a_62154_n21906# CM_p_net_0.IN a_61624_n22811# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1432 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1433 a_53562_6360# a_47184_10411# a_53040_6360# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1434 a_97830_2963# a_86263_2903# a_99787_10096# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1435 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1436 a_57294_n21906# CM_p_net_0.IN a_56456_n21906# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1437 a_50758_n27336# CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1438 a_88027_12028# a_86091_8930# PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1439 a_106442_10411# a_106442_9245# a_108378_11177# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1440 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1441 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1442 FC_top_0.AVSS a_72830_n8314# a_73230_n6322# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1443 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1444 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1445 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1446 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1447 a_n10892_n26881# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X1448 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1449 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1450 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1451 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1452 a_43602_n22894# CM_n_net_0.IN a_43042_n22894# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1453 FC_top_0.AVDD FC_top_0.IREF a_n11312_n20927# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1454 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1455 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1456 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1457 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1458 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1459 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1460 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1461 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1462 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1463 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1464 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1465 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1466 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1467 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1468 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1469 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1470 a_53194_9185# PRbiased_net_8.IBP a_60880_9245# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1471 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1472 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1473 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1474 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1475 a_62154_n36281# CM_p_net_0.IN a_61624_n39901# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1476 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1477 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1478 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1479 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1480 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1481 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1482 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1483 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1484 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1485 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1486 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1487 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1488 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1489 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1490 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1491 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1492 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1493 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1494 a_n5154_n26774# a_n11312_n21934# a_n5714_n26774# FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X1495 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1496 a_108418_n12748# a_106614_n13966# PRbiased_net_0.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1497 PRbiased_net_8.ITN a_47356_3218# a_47756_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1498 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1499 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1500 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1501 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1502 a_47714_n6773# a_47184_n7939# a_47184_n6773# PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1503 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1504 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1505 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1506 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1507 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1508 a_91947_6045# a_86091_10096# a_93873_2963# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1509 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1510 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1511 FC_top_0.VOUT a_n11312_n21934# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1512 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1513 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1514 FC_top_0.VOUT a_n11312_n21934# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1515 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1516 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1517 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1518 a_47714_n4841# a_47184_n7939# a_47184_n6773# PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1519 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1520 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1521 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1522 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1523 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1524 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1525 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1526 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1527 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1528 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1529 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1530 a_33908_n38941# CM_n_net_0.IN a_33386_n39838# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1531 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1532 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1533 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1534 a_86621_n8254# a_86091_n8254# a_86091_n8254# PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1535 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1536 a_49120_11177# a_47184_9245# PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1537 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1538 a_79110_12028# PRbiased_net_7.IBP a_72830_8870# PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1539 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1540 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1541 a_91947_2963# a_92101_8870# a_92501_8930# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1542 PRbiased_net_6.VB a_92101_8870# a_93907_8930# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1543 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1544 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1545 a_43042_n27379# CM_n_net_0.IN a_42520_n28276# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1546 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1547 a_35342_n38044# CM_n_net_0.IN a_34820_n38941# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1548 a_50758_n36281# CM_p_net_0.IN a_50228_n35376# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1549 a_120107_n12748# a_118181_n13906# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1550 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1551 a_86621_n6322# a_86091_n8254# a_86091_n8254# PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1552 a_31070_n35353# CM_n_net_0.IN a_30510_n35353# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1553 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1554 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1555 a_68796_n11139# a_66992_n14281# PRbiased_net_2.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1556 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1557 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1558 a_52164_n26431# CM_p_net_0.IN a_51596_n26431# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1559 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1560 a_49160_n11982# PRbiased_net_3.IBN PRbiased_net_3.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1561 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1562 PRbiased_net_1.ITP a_86263_n14281# a_98381_n8254# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1563 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1564 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1565 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1566 a_99787_8930# PRbiased_net_6.IBP PRbiased_net_6.ITP PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1567 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1568 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1569 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1570 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1571 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1572 a_53562_n13906# a_47184_n6773# a_53040_n13906# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1573 a_36776_n27379# CM_n_net_0.IN a_36254_n28276# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1574 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1575 a_29076_n38044# CM_n_net_0.IN a_28554_n38941# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1576 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1577 a_79081_n12297# a_78559_n14221# a_78559_n14221# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1578 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1579 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1580 a_50758_n26431# CM_p_net_0.IN a_50228_n26431# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1581 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1582 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1583 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1584 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1585 PRbiased_net_1.ITP a_86263_n14281# a_98381_n6322# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1586 a_108418_n10824# a_106614_n13966# PRbiased_net_0.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1587 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1588 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1589 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1590 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1591 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1592 a_57862_n37186# CM_p_net_0.IN a_57294_n37186# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1593 PRbiased_net_3.IBP a_53194_n7999# a_55000_n6773# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1594 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1595 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1596 a_33908_n29173# CM_n_net_0.IN a_33386_n29173# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1597 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1598 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1599 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1600 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1601 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1602 a_66820_n7088# a_66820_n8254# a_68756_n8254# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1603 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1604 a_73198_n14221# a_66820_n7088# a_72676_n14221# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1605 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1606 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1607 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1608 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1609 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1610 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1611 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1612 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1613 a_40174_n27379# CM_n_net_0.IN a_39652_n27379# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1614 a_118703_n11982# a_118181_n13906# a_118181_n13906# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1615 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1616 PRbiased_net_3.VA a_53194_n7999# a_55000_n4841# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1617 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1618 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1619 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1620 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1621 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1622 a_56456_n37186# CM_p_net_0.IN a_55926_n38091# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1623 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1624 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1625 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1626 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1627 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1628 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1629 a_66820_n7088# a_66820_n8254# a_68756_n6322# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1630 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1631 a_57862_n28241# CM_p_net_0.IN a_57294_n28241# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1632 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1633 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1634 PRbiased_net_1.VB a_92101_n8314# a_93907_n8254# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1635 a_86663_n12297# a_86263_n14281# a_86091_n8254# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1636 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1637 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1638 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1639 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1640 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1641 a_28212_9245# a_27682_9245# a_27682_9245# PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1642 a_43602_n33559# CM_n_net_0.IN a_43042_n32662# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1643 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1644 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1645 a_35902_n38044# CM_n_net_0.IN a_36776_n36250# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1646 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1647 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1648 a_120107_n10824# a_118181_n13906# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1649 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1650 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1651 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1652 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1653 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1654 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1655 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1656 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1657 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1658 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1659 PRbiased_net_1.IBP a_92101_n8314# a_93907_n6322# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1660 PRbiased_net_0.VB a_112452_n7999# a_114258_n7939# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1661 a_29658_6360# a_27854_3218# PRbiased_net_9.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1662 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1663 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1664 a_56456_n28241# CM_p_net_0.IN a_55926_n28241# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1665 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1666 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1667 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1668 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1669 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1670 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1671 a_88067_n11139# a_86263_n14281# PRbiased_net_1.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1672 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1673 PRbiased_net_4.VDD a_27682_n6773# a_35464_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1674 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1675 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1676 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1677 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1678 a_114224_6360# a_106442_10411# a_106614_3218# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1679 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1680 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1681 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1682 a_67350_10862# a_66820_8930# a_66820_8930# PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1683 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1684 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1685 a_52164_n34471# CM_p_net_0.IN a_51596_n34471# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1686 a_35902_n27379# CM_n_net_0.IN a_36776_n25585# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1687 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1688 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1689 a_52732_n27336# CM_p_net_0.IN a_52164_n27336# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1690 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1691 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1692 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1693 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1694 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1695 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1696 a_35342_n33559# CM_n_net_0.IN a_34820_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1697 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1698 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1699 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1700 a_98352_n12297# a_97830_n14221# a_97830_n14221# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1701 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1702 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1703 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1704 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1705 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1706 a_60849_4436# a_58923_3278# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1707 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1708 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1709 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1710 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1711 a_62154_n20096# CM_p_net_0.IN a_61624_n23716# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1712 a_118732_n6007# a_106614_n13966# a_118181_n13906# PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1713 a_57294_n20096# CM_p_net_0.IN a_56456_n20096# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1714 PRbiased_net_8.ITN a_47356_3218# a_47756_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1715 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1716 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1717 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1718 a_50758_n34471# CM_p_net_0.IN a_50228_n34471# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1719 a_92501_12028# a_92101_8870# PRbiased_net_6.VB PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1720 FC_top_0.AVSS a_112452_9185# a_112852_11177# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1721 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1722 a_57862_n21906# CM_p_net_0.IN a_57294_n21906# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1723 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1724 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1725 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1726 PRbiased_net_9.VDD a_27682_10411# a_35464_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1727 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1728 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1729 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1730 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1731 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1732 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1733 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1734 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1735 a_29076_n33559# CM_n_net_0.IN a_28554_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1736 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1737 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1738 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1739 a_35342_n22894# CM_n_net_0.IN a_34820_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1740 PRbiased_net_4.ITN a_27854_n13966# a_28254_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1741 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1742 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1743 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1744 PRbiased_net_4.IBN a_27682_n6773# a_34060_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1745 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1746 a_64966_n37186# CM_p_net_0.IN a_64128_n37186# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1747 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1748 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1749 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1750 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1751 a_56456_n21906# CM_p_net_0.IN a_55926_n22811# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1752 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1753 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1754 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1755 a_41378_9245# PRbiased_net_9.IBP PRbiased_net_9.ITP PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1756 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1757 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1758 FC_top_0.AVSS a_58923_n13906# a_59445_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1759 a_80485_n11139# a_78559_n14221# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1760 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1761 a_33908_n24688# CM_n_net_0.IN a_33386_n24688# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1762 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1763 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1764 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1765 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1766 a_78559_2963# a_78559_2963# a_80485_6045# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1767 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1768 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1769 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1770 a_43042_n37147# CM_n_net_0.IN a_42520_n37147# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1771 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1772 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1773 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1774 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1775 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1776 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1777 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1778 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1779 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1780 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1781 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1782 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1783 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1784 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1785 a_29076_n22894# CM_n_net_0.IN a_28554_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1786 a_5821_n12405# a_n11312_n21934# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1787 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1788 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1789 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1790 a_34060_4436# a_27682_10411# PRbiased_net_9.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1791 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1792 a_55000_n7939# a_53194_n7999# a_53040_n10824# PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1793 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1794 a_5821_n12405# a_n11312_n21934# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1795 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1796 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1797 a_72676_2963# a_72830_8870# a_73230_8930# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1798 a_33538_n13906# a_27682_n6773# a_35464_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1799 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1800 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1801 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1802 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1803 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1804 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1805 CM_p_net_0.VDD CM_p_net_0.IN a_64128_n28241# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1806 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1807 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1808 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1809 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1810 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1811 a_36776_n37147# CM_n_net_0.IN a_36254_n37147# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1812 a_56456_n36281# CM_p_net_0.IN a_55926_n39901# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1813 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1814 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1815 a_43042_n26482# CM_n_net_0.IN a_42520_n26482# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1816 PRbiased_net_7.VA a_72830_8870# a_74636_12028# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1817 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1818 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1819 a_93873_n13063# a_86091_n7088# PRbiased_net_1.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1820 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1821 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1822 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1823 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1824 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1825 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1826 a_29618_n7939# a_27682_n7939# PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1827 PRbiased_net_3.VDD a_47184_n7939# a_47714_n7939# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1828 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1829 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1830 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1831 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1832 a_79081_n14221# a_78559_n14221# a_78559_n14221# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1833 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1834 a_41608_n28276# CM_n_net_0.IN a_41086_n28276# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1835 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1836 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1837 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1838 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1839 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1840 a_n5154_n26774# a_n11312_n21934# a_n5714_n26221# FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X1841 a_40734_n36250# CM_n_net_0.IN a_40174_n36250# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1842 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1843 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1844 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1845 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1846 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1847 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1848 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1849 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1850 a_36776_n26482# CM_n_net_0.IN a_36254_n26482# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1851 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1852 a_40174_n37147# CM_n_net_0.IN a_39652_n38044# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1853 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1854 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1855 a_39972_12343# PRbiased_net_9.IBP a_33692_9185# PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1856 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1857 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1858 a_29658_n12748# a_27854_n13966# PRbiased_net_4.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1859 a_106972_n6773# a_106442_n7939# a_106442_n6773# PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1860 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1861 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1862 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1863 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1864 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1865 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1866 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1867 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1868 a_34468_n36250# CM_n_net_0.IN a_33908_n36250# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1869 a_79110_8930# a_66992_2903# a_78559_2963# PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1870 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1871 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1872 FC_top_0.AVSS a_58923_n13906# a_59445_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1873 a_40734_n25585# CM_n_net_0.IN a_40174_n25585# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1874 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1875 a_n11312_n20927# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1876 a_52732_n26431# CM_p_net_0.IN a_52164_n26431# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1877 a_39972_10411# PRbiased_net_9.IBP a_33692_9185# PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1878 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1879 a_78559_2963# a_78559_2963# a_80485_4121# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1880 a_106972_n4841# a_106442_n7939# a_106442_n6773# PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1881 a_86663_n14221# a_86263_n14281# a_86091_n8254# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1882 a_64966_n21906# CM_p_net_0.IN a_64128_n21906# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1883 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1884 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1885 a_92501_8930# a_92101_8870# PRbiased_net_6.VA PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1886 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1887 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1888 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1889 a_40174_n26482# CM_n_net_0.IN a_39652_n27379# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1890 a_33692_9185# PRbiased_net_9.IBP a_41378_11177# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1891 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1892 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1893 a_62154_n21001# CM_p_net_0.IN CM_p_net_0.OUT5 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1894 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1895 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1896 PRbiased_net_4.VDD a_27682_n7939# a_28212_n6773# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1897 a_57294_n21001# CM_p_net_0.IN a_56456_n21001# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1898 a_112820_n13906# a_106442_n6773# a_112298_n13906# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1899 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1900 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1901 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1902 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1903 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1904 a_106972_9245# a_106442_9245# a_106442_9245# PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1905 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1906 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1907 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1908 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1909 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1910 a_80516_n7088# a_66992_n14281# PRbiased_net_2.ITP PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1911 a_34468_n25585# CM_n_net_0.IN a_33908_n25585# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1912 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1913 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1914 a_58430_n37186# CM_p_net_0.IN a_57862_n37186# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1915 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1916 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1917 a_53040_3278# a_53194_9185# a_53594_9245# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1918 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1919 PRbiased_net_4.VDD a_27682_n7939# a_28212_n4841# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1920 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1921 a_37336_n35353# CM_n_net_0.IN a_36776_n35353# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1922 FC_top_0.AVSS a_92101_8870# a_92501_10862# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1923 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1924 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1925 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1926 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1927 PRbiased_net_3.VDD a_47184_n6773# a_54966_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1928 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1929 a_64966_n36281# CM_p_net_0.IN CM_p_net_0.OUT12 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1930 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1931 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1932 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1933 a_80516_n5156# a_66992_n14281# PRbiased_net_2.ITP PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1934 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1935 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1936 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1937 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1938 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1939 a_62992_n27336# CM_p_net_0.IN a_62154_n27336# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1940 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1941 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1942 FC_top_0.AVSS a_72830_n8314# a_73230_n7088# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1943 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1944 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1945 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1946 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1947 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1948 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1949 a_98352_n14221# a_97830_n14221# a_97830_n14221# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1950 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1951 a_n11312_n21934# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1952 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1953 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1954 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1955 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1956 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1957 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1958 FC_top_0.AVSS a_39421_n13906# a_39943_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1959 a_58430_n28241# CM_p_net_0.IN a_57862_n28241# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1960 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1961 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1962 a_n11312_n20927# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1963 a_29658_n10824# a_27854_n13966# PRbiased_net_4.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1964 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1965 a_72676_n11139# a_72830_n8314# a_73230_n5156# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1966 a_43042_n21997# CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1967 PRbiased_net_5.VDD a_106442_9245# a_106972_12343# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1968 FC_top_0.AVSS a_58923_3278# a_59445_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1969 a_66820_8930# a_66992_2903# a_68796_6045# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1970 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1971 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1972 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1973 a_35342_n32662# CM_n_net_0.IN a_34468_n36250# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1974 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1975 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1976 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1977 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1978 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1979 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1980 a_92101_8870# PRbiased_net_6.IBP a_99787_10862# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1981 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X1982 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1983 PRbiased_net_5.VDD a_106442_10411# a_114224_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1984 a_33908_n34456# CM_n_net_0.IN a_33386_n35353# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1985 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1986 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1987 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1988 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1989 a_39943_n11982# a_39421_n13906# a_39421_n13906# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1990 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1991 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1992 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1993 PRbiased_net_5.VDD a_106442_9245# a_106972_10411# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1994 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1995 PRbiased_net_0.IBP a_112452_n7999# a_114258_n6007# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1996 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1997 PRbiased_net_0.VDD a_106442_n6773# a_114224_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1998 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1999 a_36776_n21997# CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2000 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2001 a_29076_n32662# CM_n_net_0.IN a_28202_n36250# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2002 a_28202_n28276# CM_n_net_0.IN a_27642_n27379# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2003 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2004 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2005 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2006 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2007 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2008 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2009 a_52732_n34471# CM_p_net_0.IN a_52164_n34471# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2010 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2011 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2012 a_28212_12343# a_27682_9245# a_27682_10411# PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2013 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2014 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2015 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2016 a_n13565_n12405# a_n11312_n21934# a_5821_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2017 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2018 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2019 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2020 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2021 a_67392_6045# PRbiased_net_7.IBN a_66820_10096# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2022 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2023 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2024 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2025 a_33908_n23791# CM_n_net_0.IN a_33386_n24688# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2026 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2027 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2028 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2029 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2030 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2031 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2032 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2033 a_57862_n20096# CM_p_net_0.IN a_57294_n20096# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2034 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2035 a_28212_10411# a_27682_9245# a_27682_10411# PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2036 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2037 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2038 a_58430_n21906# CM_p_net_0.IN a_57862_n21906# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2039 a_40174_n21997# CM_n_net_0.IN a_39652_n22894# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2040 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2041 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2042 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2043 FC_top_0.AVDD FC_top_0.IREF a_n11312_n21934# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2044 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2045 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2046 a_41608_n38044# CM_n_net_0.IN a_41086_n38941# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2047 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2048 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2049 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2050 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2051 a_98381_n8254# a_86263_n14281# a_97830_n14221# PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2052 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2053 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2054 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2055 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2056 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2057 PRbiased_net_0.ITN a_106614_n13966# a_107014_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2058 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2059 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2060 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2061 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2062 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X2063 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2064 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2065 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2066 a_56456_n20096# CM_p_net_0.IN a_55926_n23716# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2067 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2068 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2069 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2070 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2071 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2072 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2073 a_66820_8930# a_66992_2903# a_68796_4121# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2074 a_86621_n7088# a_86091_n8254# a_86091_n7088# PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2075 a_98381_n6322# a_86263_n14281# a_97830_n14221# PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2076 a_30510_n28276# CM_n_net_0.IN a_29988_n28276# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2077 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2078 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2079 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2080 PRbiased_net_2.ITN PRbiased_net_2.IBN a_67392_n11139# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2081 a_114258_12343# a_112452_9185# a_112298_3278# PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2082 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2083 FC_top_0.VOUT a_n11312_n21934# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2084 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2085 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2086 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2087 a_72830_8870# a_78559_2963# a_80485_4887# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2088 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2089 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2090 a_40734_n37147# CM_n_net_0.IN a_40174_n35353# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2091 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2092 a_86621_n5156# a_86091_n8254# a_86091_n7088# PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2093 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2094 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2095 a_112298_n13906# a_106442_n6773# a_114224_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2096 a_93907_10096# a_92101_8870# FC_top_0.AVSS PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2097 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2098 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2099 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2100 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2101 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2102 a_114258_10411# a_112452_9185# FC_top_0.AVSS PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2103 PRbiased_net_1.ITP PRbiased_net_1.IBP a_98381_n7088# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2104 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2105 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2106 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2107 a_55000_n6007# a_53194_n7999# FC_top_0.AVSS PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2108 a_62992_n26431# CM_p_net_0.IN a_62154_n26431# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2109 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2110 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2111 PRbiased_net_9.VA a_33692_9185# a_35498_12343# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2112 PRbiased_net_8.ITP PRbiased_net_8.IBP a_59474_12343# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2113 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2114 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2115 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2116 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2117 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2118 a_67392_4121# PRbiased_net_7.IBN a_66820_10096# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2119 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2120 a_53194_n7999# a_58923_n13906# a_60849_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2121 FC_top_0.AVSS a_118181_n13906# a_118703_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2122 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2123 a_34468_n37147# CM_n_net_0.IN a_33908_n35353# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2124 PRbiased_net_6.VDD a_86091_8930# a_86621_10096# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2125 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2126 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2127 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2128 PRbiased_net_1.ITP PRbiased_net_1.IBP a_98381_n5156# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2129 a_29618_n6007# a_27682_n7939# PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2130 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2131 PRbiased_net_3.VDD a_47184_n7939# a_47714_n6007# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2132 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2133 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2134 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2135 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2136 a_74636_n8254# a_72830_n8314# a_72676_n11139# PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2137 PRbiased_net_9.IBP a_33692_9185# a_35498_10411# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2138 PRbiased_net_8.ITP PRbiased_net_8.IBP a_59474_10411# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2139 a_106614_3218# a_106442_10411# a_112820_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2140 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2141 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2142 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2143 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2144 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2145 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2146 a_27642_n28276# CM_n_net_0.IN a_27120_n29173# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2147 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2148 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2149 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2150 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2151 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2152 a_66820_n8254# a_66820_n8254# a_68756_n7088# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2153 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2154 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2155 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2156 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2157 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2158 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2159 a_74636_n6322# a_72830_n8314# FC_top_0.AVSS PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2160 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X2161 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2162 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2163 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2164 a_58923_3278# a_58923_3278# a_60849_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2165 a_66820_n8254# a_66820_n8254# a_68756_n5156# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2166 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2167 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2168 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2169 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2170 PRbiased_net_1.IBP a_92101_n8314# a_93907_n7088# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2171 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2172 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2173 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2174 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2175 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2176 a_64436_n23716# CM_p_net_0.IN a_64128_n20096# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2177 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2178 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2179 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2180 a_97830_2963# a_97830_2963# a_99756_6045# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2181 a_n11312_n20927# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X2182 FC_top_0.AVSS a_58923_3278# a_59445_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2183 a_72830_8870# a_78559_2963# a_80485_2963# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2184 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2185 PRbiased_net_2.VDD a_66820_n7088# a_74602_n12297# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2186 PRbiased_net_1.ITN PRbiased_net_1.IBN a_86663_n11139# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2187 a_41608_n33559# CM_n_net_0.IN a_41086_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2188 a_43602_n39838# CM_n_net_0.IN a_43042_n39838# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2189 a_57862_n21001# CM_p_net_0.IN a_57294_n21001# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2190 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2191 a_53594_9245# a_53194_9185# PRbiased_net_8.VA PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2192 a_112820_6360# a_106442_10411# a_112298_6360# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2193 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2194 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2195 a_51596_n25526# CM_p_net_0.IN a_50758_n25526# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2196 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X2197 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2198 a_53562_n12748# a_47184_n6773# PRbiased_net_3.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2199 PRbiased_net_1.VA a_92101_n8314# a_93907_n5156# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2200 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2201 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2202 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2203 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2204 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2205 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2206 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2207 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2208 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2209 a_28202_n37147# CM_n_net_0.IN a_27642_n37147# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2210 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2211 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2212 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2213 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2214 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2215 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2216 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2217 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2218 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2219 a_56456_n21001# CM_p_net_0.IN CM_p_net_0.OUT3 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2220 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2221 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2222 PRbiased_net_6.ITN PRbiased_net_6.IBN a_86663_6045# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2223 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2224 a_73198_n13063# a_66820_n7088# PRbiased_net_2.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2225 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2226 a_41608_n22894# CM_n_net_0.IN a_41086_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2227 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2228 a_112452_9185# PRbiased_net_5.IBP a_120138_9245# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2229 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2230 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2231 a_62992_n34471# CM_p_net_0.IN a_62154_n34471# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2232 a_98352_6045# a_97830_2963# a_92101_8870# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2233 a_63560_n27336# CM_p_net_0.IN a_62992_n27336# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2234 a_n11312_n20927# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2235 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2236 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2237 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2238 PRbiased_net_9.IBN a_27682_10411# a_34060_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2239 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2240 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2241 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2242 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2243 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2244 a_34060_n13906# a_27682_n6773# a_33538_n13906# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2245 a_28202_n26482# CM_n_net_0.IN a_27642_n26482# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2246 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2247 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2248 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2249 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2250 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2251 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2252 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2253 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2254 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2255 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2256 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2257 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2258 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2259 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2260 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2261 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2262 a_66820_10096# PRbiased_net_7.IBN a_68796_4887# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2263 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2264 a_30510_n38044# CM_n_net_0.IN a_29988_n38941# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2265 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2266 a_n13565_n11419# a_n11312_n21934# FC_top_0.VOUT FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2267 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2268 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2269 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2270 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2271 a_97830_2963# a_97830_2963# a_99756_4121# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2272 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2273 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2274 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2275 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2276 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2277 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2278 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2279 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2280 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2281 a_53562_n10824# a_47184_n6773# a_53040_n10824# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2282 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2283 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2284 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2285 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2286 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2287 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2288 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X2289 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2290 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2291 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2292 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2293 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2294 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2295 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2296 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2297 a_60849_3278# a_58923_3278# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2298 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2299 a_51596_n33566# CM_p_net_0.IN a_50758_n33566# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2300 a_n11312_n20927# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2301 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2302 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2303 a_80516_12028# a_66992_2903# PRbiased_net_7.ITP PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2304 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2305 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2306 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2307 a_67392_4887# a_66992_2903# a_66820_8930# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2308 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2309 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2310 PRbiased_net_6.ITN PRbiased_net_6.IBN a_86663_4121# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2311 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2312 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2313 a_58430_n20096# CM_p_net_0.IN a_57862_n20096# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2314 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2315 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2316 a_53594_n7939# a_53194_n7999# PRbiased_net_3.VA PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2317 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2318 a_42168_n27379# CM_n_net_0.IN a_41608_n27379# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2319 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2320 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2321 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2322 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2323 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2324 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2325 a_64966_n21906# CM_p_net_0.IN a_64128_n21001# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2326 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2327 a_98352_4121# a_97830_2963# a_92101_8870# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2328 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2329 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2330 FC_top_0.AVDD FC_top_0.IREF a_n11312_n21934# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2331 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2332 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2333 a_33538_6360# a_27682_10411# a_35464_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2334 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2335 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2336 a_72676_6045# a_72830_8870# a_73230_12028# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2337 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2338 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2339 a_68796_n12297# PRbiased_net_2.IBN PRbiased_net_2.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2340 a_27642_n38044# CM_n_net_0.IN a_27120_n38044# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2341 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2342 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2343 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2344 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2345 PRbiased_net_4.ITN PRbiased_net_4.IBN a_28254_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2346 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2347 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2348 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2349 a_47184_n7939# a_47184_n7939# a_49120_n6773# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2350 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2351 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2352 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2353 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2354 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2355 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2356 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2357 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2358 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2359 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2360 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2361 a_39972_11177# a_27854_3218# a_39421_3278# PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2362 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2363 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2364 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2365 a_66820_10096# PRbiased_net_7.IBN a_68796_2963# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2366 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2367 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2368 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2369 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2370 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2371 a_47184_n7939# a_47184_n7939# a_49120_n4841# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2372 PRbiased_net_9.VB a_33692_9185# a_35498_9245# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2373 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2374 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2375 a_108418_n11982# PRbiased_net_0.IBN PRbiased_net_0.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2376 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2377 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2378 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2379 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2380 a_34060_3278# a_27682_10411# a_33538_3278# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2381 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2382 PRbiased_net_0.ITP PRbiased_net_0.IBP a_118732_n6773# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2383 a_62154_n38996# CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2384 CM_n_net_0.OUT1 CM_n_net_0.IN a_27642_n21997# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2385 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2386 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2387 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2388 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2389 a_57294_n38996# CM_p_net_0.IN a_56456_n38996# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2390 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2391 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2392 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2393 a_86091_n7088# a_86091_n8254# a_88027_n8254# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2394 a_n11312_n20927# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2395 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2396 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2397 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2398 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2399 a_63560_n26431# CM_p_net_0.IN a_62992_n26431# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2400 a_47756_4436# PRbiased_net_8.IBN a_47184_10411# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2401 PRbiased_net_9.ITP PRbiased_net_9.IBP a_39972_12343# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2402 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2403 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2404 a_54966_n13906# a_47184_n6773# a_47356_n13966# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2405 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2406 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2407 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2408 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2409 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2410 a_72676_n11139# a_66820_n7088# a_74602_n14221# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2411 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2412 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2413 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2414 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2415 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2416 PRbiased_net_0.ITP PRbiased_net_0.IBP a_118732_n4841# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2417 a_86091_n7088# a_86091_n8254# a_88027_n6322# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2418 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2419 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2420 a_106442_n6773# a_106442_n7939# a_108378_n7939# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2421 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2422 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2423 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2424 a_67392_2963# a_66992_2903# a_66820_8930# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2425 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2426 a_79081_n13063# a_78559_n14221# a_72830_n8314# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2427 a_30510_n33559# CM_n_net_0.IN a_29988_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2428 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2429 PRbiased_net_9.ITP PRbiased_net_9.IBP a_39972_10411# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2430 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2431 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2432 a_41608_n32662# CM_n_net_0.IN a_40734_n36250# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2433 a_43602_n39838# CM_n_net_0.IN a_43042_n38941# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2434 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2435 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2436 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2437 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2438 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2439 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2440 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2441 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2442 a_120107_n11982# a_118181_n13906# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2443 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2444 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2445 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2446 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2447 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2448 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2449 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2450 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2451 PRbiased_net_7.ITN PRbiased_net_7.IBN a_67392_6045# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2452 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2453 PRbiased_net_4.ITN PRbiased_net_4.IBN a_28254_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2454 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2455 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2456 a_53570_n25526# CM_p_net_0.IN a_52732_n25526# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2457 a_30510_n22894# CM_n_net_0.IN a_29988_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2458 a_88067_n12297# PRbiased_net_1.IBN PRbiased_net_1.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2459 a_79081_6045# a_78559_2963# a_72830_8870# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2460 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2461 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2462 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2463 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2464 a_86663_n13063# PRbiased_net_1.IBN a_86091_n7088# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2465 a_86621_12028# a_86091_8930# a_86091_10096# PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2466 PRbiased_net_5.VDD a_106442_9245# a_106972_11177# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2467 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2468 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2469 a_51596_n32661# CM_p_net_0.IN a_50758_n32661# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2470 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2471 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2472 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2473 a_35342_n39838# CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2474 a_58430_n21001# CM_p_net_0.IN a_57862_n21001# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2475 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2476 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2477 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2478 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2479 a_112820_n12748# a_106442_n6773# PRbiased_net_0.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2480 a_92101_8870# a_97830_2963# a_99756_4887# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2481 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2482 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2483 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2484 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2485 a_27642_n33559# CM_n_net_0.IN a_27120_n33559# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2486 a_64128_n25526# CM_p_net_0.IN a_63560_n25526# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2487 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2488 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2489 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2490 a_59268_n25526# CM_p_net_0.IN a_58430_n25526# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2491 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2492 PRbiased_net_8.ITN PRbiased_net_8.IBN a_47756_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2493 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2494 a_43602_n29173# CM_n_net_0.IN a_43042_n29173# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2495 PRbiased_net_6.ITP PRbiased_net_6.IBP a_98381_12028# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2496 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2497 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2498 a_29076_n39838# CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2499 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2500 a_28212_11177# a_27682_9245# a_27682_9245# PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2501 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2502 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2503 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2504 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2505 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2506 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2507 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2508 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2509 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2510 a_63560_n34471# CM_p_net_0.IN a_62992_n34471# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2511 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2512 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2513 PRbiased_net_6.ITN a_86263_2903# a_86663_4887# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2514 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2515 FC_top_0.AVDD FC_top_0.IREF a_n11312_n20927# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2516 a_49120_n7939# a_47184_n7939# PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2517 a_27642_n22894# CM_n_net_0.IN a_27120_n22894# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2518 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2519 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2520 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2521 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2522 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2523 a_98352_n13063# a_97830_n14221# a_92101_n8314# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2524 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2525 a_60849_5202# a_58923_3278# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2526 a_98352_4887# a_97830_2963# a_97830_2963# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2527 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2528 a_80485_n12297# a_78559_n14221# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2529 FC_top_0.AVSS a_39421_n13906# a_39943_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2530 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2531 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2532 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2533 a_62154_n39901# CM_p_net_0.IN a_61624_n39901# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2534 a_66820_8930# a_66820_8930# a_68756_12028# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2535 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2536 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2537 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2538 a_57294_n39901# CM_p_net_0.IN a_56456_n39901# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2539 PRbiased_net_7.ITN PRbiased_net_7.IBN a_67392_4121# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2540 a_98381_n7088# PRbiased_net_1.IBP a_92101_n8314# PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2541 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2542 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2543 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2544 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2545 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2546 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2547 a_27682_n6773# PRbiased_net_4.IBN a_29658_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2548 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2549 PRbiased_net_9.VDD a_27682_10411# a_35464_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2550 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2551 a_31070_n27379# CM_n_net_0.IN a_30510_n27379# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2552 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2553 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2554 a_79081_4121# a_78559_2963# a_72830_8870# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2555 PRbiased_net_4.VDD a_27682_n6773# a_35464_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2556 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2557 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2558 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2559 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2560 a_112298_6360# a_106442_10411# a_114224_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2561 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2562 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2563 a_68796_n14221# PRbiased_net_2.IBN PRbiased_net_2.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2564 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2565 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2566 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2567 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2568 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2569 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2570 PRbiased_net_6.VA a_92101_8870# a_93907_12028# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2571 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2572 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2573 a_98381_n5156# PRbiased_net_1.IBP a_92101_n8314# PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2574 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2575 a_53570_n33566# CM_p_net_0.IN a_52732_n33566# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2576 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2577 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2578 a_114258_11177# a_112452_9185# FC_top_0.AVSS PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2579 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2580 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X2581 a_112820_n10824# a_106442_n6773# a_112298_n10824# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2582 a_92101_8870# a_97830_2963# a_99756_2963# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2583 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2584 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2585 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2586 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2587 a_120138_n6773# a_106614_n13966# PRbiased_net_0.ITP PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2588 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2589 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2590 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2591 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2592 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2593 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2594 a_34060_5202# a_27682_10411# PRbiased_net_9.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2595 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2596 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2597 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2598 a_64128_n33566# CM_p_net_0.IN a_63560_n33566# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2599 a_120138_n4841# a_106614_n13966# PRbiased_net_0.ITP PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2600 a_53570_n24621# CM_p_net_0.IN CM_p_net_0.OUT2 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2601 PRbiased_net_9.IBP a_33692_9185# a_35498_11177# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2602 PRbiased_net_8.ITP a_47356_3218# a_59474_11177# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2603 a_93907_10862# a_92101_8870# FC_top_0.AVSS PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2604 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2605 a_59268_n33566# CM_p_net_0.IN a_58430_n33566# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2606 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2607 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2608 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2609 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2610 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2611 a_53594_n6007# a_53194_n7999# PRbiased_net_3.IBP PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2612 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2613 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X2614 PRbiased_net_6.ITN a_86263_2903# a_86663_2963# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2615 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2616 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2617 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2618 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2619 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2620 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2621 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2622 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2623 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2624 a_98352_2963# a_97830_2963# a_97830_2963# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2625 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2626 a_74636_n7088# a_72830_n8314# FC_top_0.AVSS PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2627 FC_top_0.AVSS a_58923_n13906# a_59445_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2628 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2629 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2630 PRbiased_net_0.ITN PRbiased_net_0.IBN a_107014_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2631 FC_top_0.AVSS a_39421_n13906# a_39943_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2632 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2633 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2634 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2635 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2636 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2637 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2638 PRbiased_net_6.VDD a_86091_8930# a_86621_10862# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2639 a_43602_n24688# CM_n_net_0.IN a_43042_n24688# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2640 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2641 a_35498_9245# a_33692_9185# a_33538_6360# PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2642 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2643 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2644 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2645 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2646 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2647 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2648 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2649 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2650 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2651 a_59268_n24621# CM_p_net_0.IN CM_p_net_0.OUT4 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2652 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2653 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2654 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2655 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2656 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2657 a_74636_n5156# a_72830_n8314# a_72676_n14221# PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2658 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2659 a_30510_n32662# CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2660 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2661 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2662 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2663 FC_top_0.AVSS a_97830_2963# a_98352_6045# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2664 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2665 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2666 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2667 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2668 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2669 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2670 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2671 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2672 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2673 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2674 a_99787_10096# a_86263_2903# PRbiased_net_6.ITP PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2675 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2676 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2677 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2678 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2679 a_88067_n14221# PRbiased_net_1.IBN PRbiased_net_1.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2680 a_57862_n38996# CM_p_net_0.IN a_57294_n38996# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2681 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2682 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2683 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2684 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2685 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2686 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2687 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2688 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2689 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X2690 a_114224_n13906# a_106442_n6773# a_106614_n13966# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2691 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2692 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2693 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2694 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2695 FC_top_0.AVSS a_118181_n13906# a_118703_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2696 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2697 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2698 a_58923_n13906# a_58923_n13906# a_60849_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2699 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2700 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2701 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2702 a_112298_n13906# a_112452_n7999# a_112852_n7939# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2703 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2704 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2705 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2706 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2707 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2708 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2709 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2710 a_56456_n38996# CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2711 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2712 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2713 a_42168_n22894# CM_n_net_0.IN a_41608_n21997# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2714 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2715 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2716 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2717 a_106442_n6773# a_106442_n7939# a_108378_n6007# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2718 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2719 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2720 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2721 a_29658_n11982# PRbiased_net_4.IBN PRbiased_net_4.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2722 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2723 a_35342_n38941# CM_n_net_0.IN a_34820_n38941# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2724 a_n13565_n11419# a_n11312_n21934# FC_top_0.VOUT FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2725 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2726 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2727 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2728 a_n13565_n11419# a_n11312_n21934# FC_top_0.VOUT FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2729 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2730 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2731 a_27642_n32662# CM_n_net_0.IN a_27120_n33559# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2732 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2733 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2734 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2735 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2736 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2737 PRbiased_net_0.ITN PRbiased_net_0.IBN a_107014_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2738 a_53570_n33566# CM_p_net_0.IN a_52732_n32661# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2739 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2740 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2741 a_33692_n7999# a_39421_n13906# a_41347_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2742 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2743 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2744 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2745 a_53194_9185# a_58923_3278# a_60849_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2746 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2747 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2748 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2749 PRbiased_net_7.ITN a_66992_2903# a_67392_4887# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2750 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2751 a_29076_n38941# CM_n_net_0.IN a_28554_n38941# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2752 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2753 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2754 a_80485_n14221# a_78559_n14221# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2755 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2756 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2757 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2758 a_79081_4887# a_78559_2963# a_78559_2963# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2759 a_31070_n38044# CM_n_net_0.IN a_30510_n37147# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2760 FC_top_0.AVSS a_97830_2963# a_98352_4121# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2761 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2762 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2763 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2764 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2765 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2766 a_64128_n32661# CM_p_net_0.IN a_63560_n32661# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2767 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2768 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2769 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2770 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2771 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2772 a_59268_n33566# CM_p_net_0.IN a_58430_n32661# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2773 a_62154_n24621# CM_p_net_0.IN a_61624_n23716# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2774 PRbiased_net_5.VDD a_106442_10411# a_114224_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2775 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2776 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2777 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2778 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2779 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2780 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2781 a_35342_n29173# CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2782 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2783 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2784 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2785 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2786 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2787 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2788 a_31070_n27379# CM_n_net_0.IN a_30510_n26482# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2789 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2790 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2791 a_58923_n13906# a_58923_n13906# a_60849_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2792 FC_top_0.AVDD FC_top_0.IREF a_n11312_n20927# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2793 FC_top_0.AVSS a_118181_n13906# a_118703_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2794 a_108378_12343# a_106442_9245# PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2795 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2796 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2797 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2798 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2799 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2800 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2801 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2802 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2803 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2804 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2805 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2806 a_27854_3218# a_27682_10411# a_34060_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2807 a_88027_10096# a_86091_8930# PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2808 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2809 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2810 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2811 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2812 a_34060_n12748# a_27682_n6773# PRbiased_net_4.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2813 a_64966_n38996# CM_p_net_0.IN a_64128_n38996# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2814 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2815 a_108378_10411# a_106442_9245# PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2816 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2817 a_29076_n29173# CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2818 a_49120_n6007# a_47184_n7939# PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2819 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2820 a_62154_n38091# CM_p_net_0.IN a_61624_n38091# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2821 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2822 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2823 PRbiased_net_2.ITN a_66992_n14281# a_67392_n12297# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2824 a_57294_n38091# CM_p_net_0.IN a_56456_n38091# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2825 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2826 a_27682_9245# a_27682_9245# a_29618_12343# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2827 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2828 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2829 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2830 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2831 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2832 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2833 a_57862_n39901# CM_p_net_0.IN a_57294_n39901# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2834 a_59445_4436# a_58923_3278# a_53194_9185# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2835 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2836 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2837 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2838 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2839 a_33692_n7999# PRbiased_net_4.IBP a_41378_n7939# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2840 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2841 a_106442_n6773# PRbiased_net_0.IBN a_108418_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2842 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2843 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2844 PRbiased_net_0.VDD a_106442_n6773# a_114224_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2845 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2846 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2847 a_43602_n35353# CM_n_net_0.IN a_43042_n34456# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2848 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2849 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2850 PRbiased_net_7.ITN a_66992_2903# a_67392_2963# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2851 a_58923_3278# a_47356_3218# a_60880_12343# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2852 a_68756_n8254# a_66820_n8254# PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2853 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2854 a_27682_9245# a_27682_9245# a_29618_10411# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2855 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2856 a_79081_2963# a_78559_2963# a_78559_2963# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2857 a_56456_n39901# CM_p_net_0.IN a_55926_n39901# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2858 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2859 a_66820_n8254# a_66992_n14281# a_68796_n11139# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2860 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2861 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2862 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2863 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2864 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2865 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2866 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2867 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2868 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2869 a_58923_3278# a_47356_3218# a_60880_10411# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2870 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2871 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2872 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2873 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2874 FC_top_0.AVDD FC_top_0.IREF a_n11312_n20927# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2875 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2876 a_68756_n6322# a_66820_n8254# PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2877 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2878 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2879 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2880 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2881 a_52164_n37186# CM_p_net_0.IN a_51596_n37186# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2882 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2883 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2884 a_47356_n13966# a_47184_n6773# a_53562_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2885 a_43602_n24688# CM_n_net_0.IN a_43042_n23791# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2886 a_37336_n27379# CM_n_net_0.IN a_36776_n27379# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2887 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2888 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2889 FC_top_0.AVSS a_78559_2963# a_79081_6045# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2890 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2891 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2892 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2893 a_86091_n8254# a_86091_n8254# a_88027_n7088# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2894 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2895 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2896 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2897 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2898 PRbiased_net_9.ITP a_27854_3218# a_39972_11177# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2899 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2900 a_62154_n31756# CM_p_net_0.IN a_61624_n35376# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2901 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2902 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2903 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2904 a_57294_n31756# CM_p_net_0.IN a_56456_n31756# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2905 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2906 a_50758_n37186# CM_p_net_0.IN a_50228_n38091# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2907 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2908 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2909 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2910 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2911 a_86091_n8254# a_86091_n8254# a_88027_n5156# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2912 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2913 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2914 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2915 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2916 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2917 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2918 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2919 a_112852_9245# a_112452_9185# PRbiased_net_5.VA PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2920 a_34060_n10824# a_27682_n6773# a_33538_n10824# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2921 a_52164_n28241# CM_p_net_0.IN a_51596_n28241# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2922 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2923 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2924 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2925 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2926 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2927 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2928 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2929 a_79110_10096# PRbiased_net_7.IBP a_72830_8870# PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2930 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2931 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2932 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2933 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2934 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2935 a_41608_n39838# CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2936 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2937 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2938 FC_top_0.AVSS a_58923_3278# a_59445_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2939 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2940 PRbiased_net_1.ITN a_86263_n14281# a_86663_n12297# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2941 a_31070_n22894# CM_n_net_0.IN a_30510_n21997# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2942 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2943 a_62154_n22811# CM_p_net_0.IN a_61624_n22811# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2944 a_98381_12028# PRbiased_net_6.IBP a_92101_8870# PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2945 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2946 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2947 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2948 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2949 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2950 a_57294_n22811# CM_p_net_0.IN a_56456_n22811# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2951 a_50758_n28241# CM_p_net_0.IN a_50228_n28241# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2952 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2953 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2954 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2955 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2956 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2957 a_53194_9185# a_58923_3278# a_60849_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2958 FC_top_0.AVSS a_97830_2963# a_98352_4887# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2959 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2960 a_58430_n38996# CM_p_net_0.IN a_57862_n38996# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2961 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2962 a_n5714_n27397# a_n11312_n21934# a_n6236_n27397# FC_top_0.AVSS nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X2963 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2964 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2965 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2966 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2967 a_47756_3278# a_47356_3218# a_47184_9245# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2968 CM_p_net_0.VDD CM_p_net_0.IN a_64128_n39901# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2969 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2970 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2971 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2972 a_54966_n12748# a_47184_n6773# PRbiased_net_3.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2973 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2974 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2975 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2976 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2977 PRbiased_net_2.VDD a_66820_n7088# a_74602_n13063# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2978 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2979 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2980 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2981 FC_top_0.AVSS a_78559_2963# a_79081_4121# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2982 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2983 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2984 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2985 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2986 a_n11312_n20927# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2987 a_43042_n28276# CM_n_net_0.IN a_42520_n28276# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2988 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2989 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2990 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2991 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2992 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2993 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2994 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2995 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2996 FC_top_0.AVSS a_112452_n7999# a_112852_n6007# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2997 a_52164_n21906# CM_p_net_0.IN a_51596_n21906# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2998 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2999 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3000 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3001 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3002 a_34092_n6773# a_33692_n7999# PRbiased_net_4.IBP PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3003 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3004 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3005 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3006 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3007 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3008 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3009 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3010 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3011 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3012 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3013 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3014 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3015 a_36776_n28276# CM_n_net_0.IN a_36254_n28276# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3016 a_50758_n21906# CM_p_net_0.IN a_50228_n22811# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3017 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3018 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3019 a_112452_n7999# a_118181_n13906# a_120107_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3020 PRbiased_net_9.IBN a_27682_10411# a_34060_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3021 a_74636_12028# a_72830_8870# a_72676_2963# PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3022 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3023 a_34092_n4841# a_33692_n7999# PRbiased_net_4.VB PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3024 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3025 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3026 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3027 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3028 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3029 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3030 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3031 a_47756_n13906# a_47356_n13966# a_47184_n7939# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3032 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3033 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3034 a_98381_8930# a_86263_2903# a_97830_2963# PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3035 a_53562_n11982# a_47184_n6773# PRbiased_net_3.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3036 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3037 PRbiased_net_2.ITN a_66992_n14281# a_67392_n14221# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3038 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3039 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3040 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3041 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3042 a_40734_n28276# CM_n_net_0.IN a_40174_n27379# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3043 a_78559_n14221# a_78559_n14221# a_80485_n11139# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3044 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3045 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3046 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3047 a_40174_n28276# CM_n_net_0.IN a_39652_n29173# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3048 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3049 FC_top_0.AVSS a_97830_2963# a_98352_2963# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3050 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3051 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3052 a_66820_10096# a_66820_8930# a_68756_8930# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3053 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3054 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3055 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3056 a_n11312_n20927# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3057 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3058 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3059 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3060 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3061 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3062 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3063 a_50758_n36281# CM_p_net_0.IN a_50228_n39901# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3064 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3065 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3066 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3067 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3068 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3069 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3070 a_54966_n10824# a_47184_n6773# a_47356_n13966# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3071 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3072 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3073 a_34468_n28276# CM_n_net_0.IN a_33908_n27379# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3074 a_112852_12343# a_112452_9185# PRbiased_net_5.VB PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3075 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3076 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3077 a_37336_n38044# CM_n_net_0.IN a_36776_n37147# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3078 a_120107_4436# a_118181_3278# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3079 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3080 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3081 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3082 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3083 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3084 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3085 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3086 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3087 a_92501_10096# a_92101_8870# PRbiased_net_6.IBP PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3088 a_56456_n24621# CM_p_net_0.IN a_55926_n23716# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3089 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3090 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3091 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3092 a_88027_8930# a_86091_8930# PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3093 a_112852_10411# a_112452_9185# PRbiased_net_5.IBP PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3094 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3095 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3096 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3097 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3098 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3099 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3100 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3101 a_57862_n38091# CM_p_net_0.IN a_57294_n38091# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3102 a_33538_6360# a_33692_9185# a_34092_12343# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3103 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3104 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3105 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3106 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3107 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3108 a_58430_n39901# CM_p_net_0.IN a_57862_n39901# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3109 a_118181_n13906# a_106614_n13966# a_120138_n6773# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3110 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3111 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3112 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3113 a_107014_4436# PRbiased_net_5.IBN a_106442_10411# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3114 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3115 a_37336_n27379# CM_n_net_0.IN a_36776_n26482# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3116 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3117 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3118 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3119 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3120 a_27682_n7939# a_27854_n13966# a_29658_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3121 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3122 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3123 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3124 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3125 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3126 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3127 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3128 a_35342_n34456# CM_n_net_0.IN a_34820_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3129 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3130 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3131 FC_top_0.AVSS a_33692_9185# a_34092_10411# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3132 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3133 a_33692_n7999# PRbiased_net_4.IBP a_41378_n6007# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3134 a_68796_n13063# a_66992_n14281# PRbiased_net_2.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3135 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3136 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3137 a_56456_n38091# CM_p_net_0.IN a_55926_n38091# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3138 FC_top_0.AVDD FC_top_0.IREF a_n11312_n21934# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3139 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3140 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3141 a_118181_n13906# a_106614_n13966# a_120138_n4841# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3142 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3143 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3144 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3145 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3146 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3147 a_92469_n11139# a_86091_n7088# a_91947_n11139# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3148 a_33908_n36250# CM_n_net_0.IN CM_n_net_0.OUT10 FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3149 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3150 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3151 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3152 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3153 PRbiased_net_1.ITN a_86263_n14281# a_86663_n14221# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3154 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3155 a_30510_n39838# CM_n_net_0.IN a_28202_n39838# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3156 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3157 a_52732_n37186# CM_p_net_0.IN a_52164_n37186# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3158 a_29076_n34456# CM_n_net_0.IN a_28554_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3159 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3160 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3161 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3162 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3163 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3164 a_41608_n38941# CM_n_net_0.IN a_41086_n38941# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3165 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3166 a_35342_n23791# CM_n_net_0.IN a_34820_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3167 PRbiased_net_7.IBP a_72830_8870# a_74636_10096# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3168 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3169 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3170 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3171 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3172 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3173 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3174 a_99787_10862# PRbiased_net_6.IBP PRbiased_net_6.ITP PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3175 a_88067_6045# a_86263_2903# PRbiased_net_6.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3176 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3177 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3178 FC_top_0.AVSS a_78559_2963# a_79081_4887# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3179 a_33908_n25585# CM_n_net_0.IN CM_n_net_0.OUT4 FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3180 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3181 a_47756_5202# a_47356_3218# a_47184_9245# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3182 a_43042_n38044# CM_n_net_0.IN a_42520_n38941# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3183 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3184 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3185 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3186 a_57862_n31756# CM_p_net_0.IN a_57294_n31756# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3187 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3188 a_n10892_n26881# a_n10892_n26881# a_n540_n21552# FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.78p ps=3.7u w=1.2u l=2u
X3189 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3190 PRbiased_net_4.ITN a_27854_n13966# a_28254_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3191 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3192 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3193 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3194 a_35464_4436# a_27682_10411# PRbiased_net_9.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3195 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3196 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3197 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3198 a_52732_n28241# CM_p_net_0.IN a_52164_n28241# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3199 a_29076_n23791# CM_n_net_0.IN a_28554_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3200 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3201 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3202 PRbiased_net_6.ITP a_86263_2903# a_98381_8930# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3203 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3204 a_64966_n24621# CM_p_net_0.IN a_64436_n23716# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3205 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3206 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3207 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3208 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3209 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3210 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3211 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3212 a_56456_n31756# CM_p_net_0.IN a_55926_n35376# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3213 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3214 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3215 a_41378_12343# a_27854_3218# PRbiased_net_9.ITP PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3216 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3217 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3218 a_36776_n38044# CM_n_net_0.IN a_36254_n38941# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3219 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3220 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3221 a_80485_6045# a_78559_2963# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3222 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3223 a_27682_n7939# a_27854_n13966# a_29658_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3224 a_27642_n39838# CM_n_net_0.IN a_27120_n39838# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3225 a_57862_n22811# CM_p_net_0.IN a_57294_n22811# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3226 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3227 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3228 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3229 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3230 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3231 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3232 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3233 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3234 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3235 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3236 a_41608_n29173# CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3237 a_41378_10411# a_27854_3218# PRbiased_net_9.ITP PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3238 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3239 a_88067_n13063# a_86263_n14281# PRbiased_net_1.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3240 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3241 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3242 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3243 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3244 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3245 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3246 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3247 a_40734_n37147# CM_n_net_0.IN a_40174_n37147# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3248 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3249 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3250 a_64966_n38996# CM_p_net_0.IN a_64128_n38091# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3251 FC_top_0.AVSS a_53194_n7999# a_53594_n6773# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3252 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3253 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3254 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3255 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3256 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3257 a_56456_n22811# CM_p_net_0.IN a_55926_n22811# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3258 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3259 a_40174_n38044# CM_n_net_0.IN a_39652_n38044# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3260 a_114224_n12748# a_106442_n6773# PRbiased_net_0.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3261 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3262 a_37336_n22894# CM_n_net_0.IN a_36776_n21997# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3263 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3264 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3265 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3266 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3267 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3268 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3269 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3270 a_52164_n20096# CM_p_net_0.IN a_51596_n20096# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3271 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3272 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3273 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3274 a_60849_6360# a_58923_3278# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3275 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3276 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3277 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3278 a_53040_n10824# a_53194_n7999# a_53594_n4841# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3279 a_52732_n21906# CM_p_net_0.IN a_52164_n21906# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3280 a_86091_8930# a_86091_8930# a_88027_12028# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3281 a_88067_4121# a_86263_2903# PRbiased_net_6.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3282 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3283 a_34468_n37147# CM_n_net_0.IN a_33908_n37147# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3284 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3285 FC_top_0.AVSS a_78559_2963# a_79081_2963# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3286 a_40734_n26482# CM_n_net_0.IN a_40174_n26482# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3287 a_60880_12343# a_47356_3218# PRbiased_net_8.ITP PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3288 a_108378_11177# a_106442_9245# PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3289 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3290 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3291 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3292 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3293 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3294 a_33538_3278# a_27682_10411# a_35464_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3295 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3296 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3297 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3298 a_50758_n20096# CM_p_net_0.IN a_50228_n23716# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3299 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3300 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3301 a_39972_n7939# a_27854_n13966# a_39421_n13906# PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3302 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3303 a_60880_10411# a_47356_3218# PRbiased_net_8.ITP PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3304 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3305 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3306 a_39421_n13906# a_39421_n13906# a_41347_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3307 a_35498_12343# a_33692_9185# a_33538_3278# PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3308 a_59474_12343# PRbiased_net_8.IBP a_53194_9185# PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3309 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3310 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3311 a_34468_n26482# CM_n_net_0.IN a_33908_n26482# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3312 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3313 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3314 a_107014_n13906# a_106614_n13966# a_106442_n7939# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3315 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3316 a_80485_4121# a_78559_2963# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3317 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3318 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3319 a_80485_n13063# a_78559_n14221# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3320 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3321 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X3322 a_27682_10411# a_27682_9245# a_29618_11177# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3323 a_68756_8930# a_66820_8930# PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3324 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3325 a_88027_10862# a_86091_8930# PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3326 a_112820_n11982# a_106442_n6773# PRbiased_net_0.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3327 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3328 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3329 a_64436_n35376# CM_p_net_0.IN a_64128_n31756# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3330 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3331 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3332 a_43042_n33559# CM_n_net_0.IN a_42520_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3333 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3334 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3335 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3336 a_5821_n12405# a_n11312_n21934# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3337 a_35498_10411# a_33692_9185# FC_top_0.AVSS PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3338 a_59474_10411# PRbiased_net_8.IBP a_53194_9185# PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3339 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3340 a_5821_n12405# a_n11312_n21934# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3341 a_53194_9185# PRbiased_net_8.IBP a_60880_11177# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3342 a_34060_6360# a_27682_10411# a_33538_6360# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3343 a_49160_4436# a_47356_3218# PRbiased_net_8.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3344 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3345 a_68756_n7088# a_66820_n8254# PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3346 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3347 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3348 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3349 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3350 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3351 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3352 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3353 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3354 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3355 FC_top_0.AVSS a_n11312_n20927# a_n10892_n26881# FC_top_0.AVSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X3356 a_114224_n10824# a_106442_n6773# a_106614_n13966# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3357 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3358 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3359 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3360 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3361 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3362 a_36776_n33559# CM_n_net_0.IN a_36254_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3363 a_43042_n22894# CM_n_net_0.IN a_42520_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3364 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3365 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3366 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3367 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3368 a_68756_n5156# a_66820_n8254# PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3369 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3370 a_64966_n25526# CM_p_net_0.IN a_64128_n22811# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3371 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3372 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3373 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3374 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3375 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3376 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3377 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3378 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3379 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3380 FC_top_0.AVSS a_39421_n13906# a_39943_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3381 a_62992_n37186# CM_p_net_0.IN a_62154_n37186# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3382 a_33692_9185# PRbiased_net_9.IBP a_41378_9245# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3383 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3384 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3385 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3386 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3387 a_33908_n35353# CM_n_net_0.IN a_33386_n35353# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3388 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3389 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3390 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3391 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3392 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3393 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3394 a_58430_n38091# CM_p_net_0.IN a_57862_n38091# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3395 a_30510_n38941# CM_n_net_0.IN a_29988_n38941# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3396 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3397 a_36776_n22894# CM_n_net_0.IN a_36254_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3398 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3399 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3400 a_40174_n33559# CM_n_net_0.IN a_39652_n33559# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3401 a_28202_n28276# CM_n_net_0.IN a_27642_n28276# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3402 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3403 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3404 a_59445_3278# a_58923_3278# a_58923_3278# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3405 a_68796_6045# a_66992_2903# PRbiased_net_7.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3406 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3407 PRbiased_net_0.VDD a_106442_n7939# a_106972_n7939# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3408 a_106442_n7939# a_106614_n13966# a_108418_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3409 a_39421_n13906# a_39421_n13906# a_41347_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3410 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X3411 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3412 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3413 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3414 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3415 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3416 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3417 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3418 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3419 a_62992_n28241# CM_p_net_0.IN a_62154_n28241# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3420 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3421 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3422 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3423 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3424 CM_n_net_0.OUT5 CM_n_net_0.IN a_40174_n21997# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3425 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3426 a_52164_n21001# CM_p_net_0.IN a_51596_n21001# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3427 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3428 a_n13565_n11419# a_n11312_n21934# FC_top_0.VOUT FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3429 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3430 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X3431 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3432 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3433 PRbiased_net_7.ITP a_66992_2903# a_79110_8930# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3434 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3435 a_40174_n22894# CM_n_net_0.IN a_39652_n22894# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3436 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3437 a_79110_10862# a_66992_2903# a_78559_2963# PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3438 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3439 a_49120_9245# a_47184_9245# PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3440 FC_top_0.VOUT a_n11312_n21934# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3441 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3442 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3443 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3444 FC_top_0.VOUT a_n11312_n21934# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3445 a_28212_n7939# a_27682_n7939# a_27682_n7939# PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3446 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3447 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3448 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3449 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3450 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3451 PRbiased_net_3.IBN a_47184_n6773# a_53562_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3452 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3453 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3454 a_50758_n21001# CM_p_net_0.IN CM_p_net_0.OUT1 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3455 a_47714_12343# a_47184_9245# a_47184_10411# PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3456 CM_n_net_0.OUT3 CM_n_net_0.IN a_33908_n21997# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3457 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3458 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3459 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3460 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3461 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3462 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3463 a_27642_n38941# CM_n_net_0.IN a_27120_n39838# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3464 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3465 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3466 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3467 a_30510_n29173# CM_n_net_0.IN a_28202_n29173# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3468 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3469 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3470 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3471 a_58430_n31756# CM_p_net_0.IN a_57862_n31756# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3472 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3473 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3474 PRbiased_net_0.ITN a_106614_n13966# a_107014_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3475 a_88067_4887# PRbiased_net_6.IBN PRbiased_net_6.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3476 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3477 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3478 a_47714_10411# a_47184_9245# a_47184_10411# PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3479 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3480 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3481 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3482 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3483 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3484 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3485 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3486 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3487 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3488 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3489 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3490 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3491 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3492 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3493 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3494 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3495 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3496 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3497 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3498 a_62992_n21906# CM_p_net_0.IN a_62154_n21906# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3499 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3500 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3501 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3502 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3503 FC_top_0.AVSS a_118181_3278# a_118703_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3504 a_51596_n27336# CM_p_net_0.IN a_50758_n27336# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3505 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3506 PRbiased_net_5.VDD a_106442_9245# a_106972_9245# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3507 a_68796_4121# a_66992_2903# PRbiased_net_7.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3508 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3509 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3510 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3511 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3512 a_106442_n7939# a_106614_n13966# a_108418_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3513 a_58430_n22811# CM_p_net_0.IN a_57862_n22811# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3514 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3515 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3516 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3517 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3518 a_114258_n7939# a_112452_n7999# a_112298_n10824# PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3519 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3520 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3521 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3522 a_80485_4887# a_78559_2963# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3523 a_112298_3278# a_106442_10411# a_114224_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3524 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3525 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3526 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3527 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3528 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3529 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3530 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3531 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3532 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3533 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3534 a_53194_n7999# a_58923_n13906# a_60849_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3535 a_27642_n29173# CM_n_net_0.IN a_27120_n29173# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3536 FC_top_0.AVSS a_118181_n13906# a_118703_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3537 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3538 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3539 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3540 a_n540_n22863# a_n10892_n26881# a_n1108_n22277# FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X3541 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3542 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3543 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3544 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3545 PRbiased_net_8.ITP a_47356_3218# a_59474_9245# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3546 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3547 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3548 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3549 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3550 PRbiased_net_4.VB a_33692_n7999# a_35498_n7939# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3551 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3552 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3553 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3554 PRbiased_net_3.ITP a_47356_n13966# a_59474_n7939# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3555 a_47356_n13966# a_47184_n6773# a_53562_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3556 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3557 a_118703_4436# a_118181_3278# a_112452_9185# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3558 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3559 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3560 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3561 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3562 a_52732_n20096# CM_p_net_0.IN a_52164_n20096# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3563 PRbiased_net_8.VA a_53194_9185# a_55000_12343# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3564 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3565 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3566 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3567 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3568 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3569 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3570 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3571 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3572 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3573 a_43042_n32662# CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3574 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3575 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3576 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3577 a_112852_11177# a_112452_9185# PRbiased_net_5.IBP PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3578 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3579 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3580 a_88067_2963# PRbiased_net_6.IBN PRbiased_net_6.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3581 PRbiased_net_8.IBP a_53194_9185# a_55000_10411# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3582 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3583 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3584 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3585 a_118732_n6773# PRbiased_net_0.IBP a_112452_n7999# PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3586 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3587 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3588 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3589 a_41608_n34456# CM_n_net_0.IN a_41086_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3590 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3591 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3592 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3593 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3594 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3595 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3596 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3597 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3598 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3599 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3600 a_118181_n13906# a_118181_n13906# a_120107_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3601 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3602 a_35902_n27379# CM_n_net_0.IN a_35342_n27379# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3603 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3604 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3605 a_39972_n6007# a_27854_n13966# a_39421_n13906# PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3606 a_36776_n32662# CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3607 a_28202_n38941# CM_n_net_0.IN a_27642_n38044# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3608 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3609 a_66820_n7088# PRbiased_net_2.IBN a_68796_n12297# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3610 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3611 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3612 FC_top_0.AVSS a_33692_9185# a_34092_11177# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3613 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3614 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3615 a_86091_8930# a_86263_2903# a_88067_6045# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3616 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3617 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3618 a_118732_n4841# PRbiased_net_0.IBP a_112452_n7999# PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3619 a_92501_10862# a_92101_8870# PRbiased_net_6.IBP PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3620 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3621 a_47756_n12748# PRbiased_net_3.IBN a_47184_n6773# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3622 a_30510_n24688# CM_n_net_0.IN a_29988_n26482# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3623 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3624 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3625 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3626 a_41347_4436# a_39421_3278# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3627 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3628 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3629 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3630 PRbiased_net_2.ITN PRbiased_net_2.IBN a_67392_n13063# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3631 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3632 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3633 a_99756_6045# a_97830_2963# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3634 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3635 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3636 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3637 a_41608_n23791# CM_n_net_0.IN a_41086_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3638 a_59445_5202# a_58923_3278# a_58923_3278# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3639 a_73198_6045# a_66820_10096# a_72676_6045# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3640 a_80485_2963# a_78559_2963# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3641 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X3642 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3643 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3644 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3645 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3646 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3647 a_29636_n27379# CM_n_net_0.IN a_29076_n27379# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3648 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3649 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3650 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3651 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3652 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3653 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3654 a_40174_n32662# CM_n_net_0.IN a_39652_n33559# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3655 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3656 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3657 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3658 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3659 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3660 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3661 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3662 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3663 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3664 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3665 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3666 a_80516_10096# a_66992_2903# PRbiased_net_7.ITP PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3667 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3668 a_86663_6045# PRbiased_net_6.IBN a_86091_10096# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3669 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3670 a_120107_3278# a_118181_3278# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3671 a_28254_n13906# a_27854_n13966# a_27682_n7939# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3672 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3673 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3674 a_34060_n11982# a_27682_n6773# PRbiased_net_4.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3675 a_51596_n26431# CM_p_net_0.IN a_50758_n26431# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3676 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3677 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3678 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3679 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3680 a_63560_n37186# CM_p_net_0.IN a_62992_n37186# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3681 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3682 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3683 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3684 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3685 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3686 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3687 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3688 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3689 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3690 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3691 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3692 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3693 a_27642_n24688# CM_n_net_0.IN a_27120_n24688# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3694 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3695 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3696 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3697 a_n540_n21552# a_n10892_n26881# a_n1108_n21552# FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X3698 PRbiased_net_7.IBP a_72830_8870# a_74636_10862# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3699 FC_top_0.AVSS a_72830_8870# a_73230_10096# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3700 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3701 a_n13565_n12405# a_n11312_n21934# a_5821_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3702 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3703 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3704 a_107014_3278# a_106614_3218# a_106442_9245# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3705 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3706 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3707 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3708 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3709 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3710 a_118181_n13906# a_118181_n13906# a_120107_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3711 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3712 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3713 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3714 a_5821_n12405# a_n11312_n21934# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3715 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3716 a_58923_3278# a_58923_3278# a_60849_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3717 a_63560_n28241# CM_p_net_0.IN a_62992_n28241# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3718 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3719 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3720 a_5821_n12405# a_n11312_n21934# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3721 a_68796_4887# PRbiased_net_7.IBN PRbiased_net_7.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3722 a_86091_8930# a_86263_2903# a_88067_4121# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3723 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3724 PRbiased_net_0.VDD a_106442_n7939# a_106972_n6007# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3725 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3726 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3727 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3728 a_47756_n10824# PRbiased_net_3.IBN a_47184_n6773# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3729 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3730 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3731 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3732 a_52732_n21001# CM_p_net_0.IN a_52164_n21001# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3733 a_41378_11177# PRbiased_net_9.IBP PRbiased_net_9.ITP PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3734 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3735 a_99756_4121# a_97830_2963# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3736 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3737 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3738 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3739 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3740 a_42168_n29173# CM_n_net_0.IN a_41608_n28276# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3741 a_73198_4121# a_66820_10096# PRbiased_net_7.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3742 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3743 PRbiased_net_1.ITN PRbiased_net_1.IBN a_86663_n13063# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3744 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3745 a_n1108_n22277# a_n10892_n26881# a_n1676_n22277# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X3746 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3747 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3748 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3749 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3750 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3751 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3752 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3753 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3754 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3755 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3756 a_68756_12028# a_66820_8930# PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3757 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3758 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3759 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3760 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3761 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3762 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3763 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3764 a_28212_n6007# a_27682_n7939# a_27682_n7939# PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3765 a_28202_n34456# CM_n_net_0.IN a_27642_n33559# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3766 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3767 a_73230_n8254# a_72830_n8314# PRbiased_net_2.VA PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3768 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3769 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3770 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3771 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3772 a_86663_4121# PRbiased_net_6.IBN a_86091_10096# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3773 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3774 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3775 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3776 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3777 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3778 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3779 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3780 a_53570_n27336# CM_p_net_0.IN a_52732_n27336# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3781 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3782 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3783 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3784 a_27854_3218# a_27682_10411# a_34060_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3785 a_35464_3278# a_27682_10411# a_27854_3218# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3786 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3787 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3788 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3789 a_47184_9245# a_47356_3218# a_49160_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3790 a_73230_n6322# a_72830_n8314# PRbiased_net_2.IBP PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3791 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3792 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3793 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3794 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3795 a_62992_n20096# CM_p_net_0.IN a_62154_n20096# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3796 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3797 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3798 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3799 a_28202_n23791# CM_n_net_0.IN a_27642_n22894# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3800 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3801 a_60880_11177# PRbiased_net_8.IBP PRbiased_net_8.ITP PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3802 a_63560_n21906# CM_p_net_0.IN a_62992_n21906# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3803 a_106614_n13966# a_106442_n6773# a_112820_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3804 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3805 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3806 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3807 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3808 a_51596_n34471# CM_p_net_0.IN a_50758_n34471# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3809 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3810 a_106972_12343# a_106442_9245# a_106442_10411# PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3811 a_47184_n6773# PRbiased_net_3.IBN a_49160_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3812 a_72830_n8314# a_78559_n14221# a_80485_n12297# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3813 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3814 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3815 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3816 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3817 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3818 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3819 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3820 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3821 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3822 a_64128_n27336# CM_p_net_0.IN a_63560_n27336# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3823 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3824 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3825 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3826 a_59268_n27336# CM_p_net_0.IN a_58430_n27336# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3827 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3828 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3829 a_68796_2963# PRbiased_net_7.IBN PRbiased_net_7.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3830 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3831 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3832 a_86621_10096# a_86091_8930# a_86091_10096# PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3833 a_35498_11177# a_33692_9185# FC_top_0.AVSS PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3834 a_59474_11177# a_47356_3218# a_58923_3278# PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3835 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3836 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3837 a_59474_9245# a_47356_3218# a_58923_3278# PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3838 a_106972_10411# a_106442_9245# a_106442_10411# PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3839 a_30510_n34456# CM_n_net_0.IN a_29988_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3840 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3841 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3842 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3843 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3844 a_114258_n6007# a_112452_n7999# FC_top_0.AVSS PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3845 a_54966_n11982# a_47184_n6773# PRbiased_net_3.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3846 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3847 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3848 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3849 a_66820_n7088# PRbiased_net_2.IBN a_68796_n14221# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3850 PRbiased_net_9.VDD a_27682_9245# a_28212_12343# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3851 a_86263_2903# a_86091_10096# a_92469_6045# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3852 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3853 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3854 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3855 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3856 PRbiased_net_0.IBP a_112452_n7999# a_114258_n6773# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3857 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3858 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3859 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3860 PRbiased_net_4.ITP a_27854_n13966# a_39972_n7939# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3861 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3862 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3863 FC_top_0.AVDD FC_top_0.IREF a_n11312_n21934# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3864 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3865 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3866 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3867 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3868 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3869 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3870 PRbiased_net_6.ITP PRbiased_net_6.IBP a_98381_10096# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3871 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3872 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3873 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3874 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3875 PRbiased_net_9.VDD a_27682_9245# a_28212_10411# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3876 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3877 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3878 PRbiased_net_4.IBP a_33692_n7999# a_35498_n6007# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3879 PRbiased_net_3.ITP a_47356_n13966# a_59474_n6007# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3880 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3881 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3882 a_30510_n23791# CM_n_net_0.IN a_29988_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3883 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3884 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3885 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3886 a_72830_n8314# PRbiased_net_2.IBP a_80516_n8254# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3887 PRbiased_net_0.VA a_112452_n7999# a_114258_n4841# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3888 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3889 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3890 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3891 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3892 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X3893 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3894 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3895 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3896 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3897 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3898 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3899 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3900 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3901 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3902 a_n1108_n21552# a_n10892_n26881# a_n1676_n21552# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X3903 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3904 a_120107_5202# a_118181_3278# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3905 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3906 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3907 a_72830_n8314# PRbiased_net_2.IBP a_80516_n6322# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3908 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3909 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3910 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3911 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3912 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3913 PRbiased_net_2.ITP a_66992_n14281# a_79110_n8254# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3914 a_66820_8930# a_66820_8930# a_68756_10096# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3915 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3916 a_53570_n36281# CM_p_net_0.IN a_53040_n35376# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3917 a_27642_n34456# CM_n_net_0.IN a_27120_n35353# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3918 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3919 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3920 a_92469_n12297# a_86091_n7088# PRbiased_net_1.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3921 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3922 a_107014_n12748# PRbiased_net_0.IBN a_106442_n6773# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3923 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3924 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3925 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3926 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3927 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3928 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3929 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3930 PRbiased_net_2.ITP a_66992_n14281# a_79110_n6322# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3931 a_91947_n14221# a_86091_n7088# a_93873_n11139# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3932 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3933 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3934 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3935 a_86091_10096# PRbiased_net_6.IBN a_88067_4887# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3936 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3937 PRbiased_net_6.IBP a_92101_8870# a_93907_10096# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3938 a_107014_5202# a_106614_3218# a_106442_9245# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3939 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3940 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3941 a_52164_n38996# CM_p_net_0.IN a_51596_n38996# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3942 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3943 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3944 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3945 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3946 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3947 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3948 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3949 a_49160_3278# PRbiased_net_8.IBN PRbiased_net_8.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3950 a_99756_4887# a_97830_2963# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3951 a_27642_n23791# CM_n_net_0.IN a_27120_n24688# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3952 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3953 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3954 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3955 a_53570_n27336# CM_p_net_0.IN a_52732_n26431# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3956 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3957 a_73198_4887# a_66820_10096# PRbiased_net_7.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3958 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3959 a_42168_n38044# CM_n_net_0.IN a_41608_n38044# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3960 a_59268_n36281# CM_p_net_0.IN a_58738_n35376# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3961 PRbiased_net_6.IBN a_86091_10096# a_92469_4121# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3962 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3963 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3964 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3965 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3966 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3967 a_47756_6360# PRbiased_net_8.IBN a_47184_10411# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3968 FC_top_0.AVDD a_n10892_n26881# a_n1108_n23588# FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X3969 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3970 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3971 a_62992_n21001# CM_p_net_0.IN a_62154_n21001# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3972 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3973 a_55000_n6773# a_53194_n7999# FC_top_0.AVSS PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3974 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3975 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3976 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3977 a_50758_n38996# CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3978 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3979 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3980 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3981 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3982 a_31070_n29173# CM_n_net_0.IN a_30510_n28276# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3983 FC_top_0.AVDD FC_top_0.IREF a_n11312_n20927# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3984 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3985 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3986 a_86663_4887# a_86263_2903# a_86091_8930# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3987 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3988 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3989 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3990 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3991 a_47714_11177# a_47184_9245# a_47184_9245# PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3992 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3993 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3994 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3995 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3996 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3997 a_64128_n26431# CM_p_net_0.IN a_63560_n26431# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3998 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3999 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4000 a_55000_n4841# a_53194_n7999# a_53040_n13906# PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4001 a_67392_n11139# PRbiased_net_2.IBN a_66820_n7088# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4002 a_59268_n27336# CM_p_net_0.IN a_58430_n26431# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4003 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4004 a_29618_n6773# a_27682_n7939# PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4005 PRbiased_net_3.VDD a_47184_n7939# a_47714_n6773# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4006 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4007 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4008 a_27682_n6773# PRbiased_net_4.IBN a_29658_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4009 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4010 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4011 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4012 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4013 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4014 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4015 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4016 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4017 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4018 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4019 a_35902_n22894# CM_n_net_0.IN a_35342_n21997# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4020 FC_top_0.VOUT a_n11312_n21934# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4021 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4022 CM_n_net_0.OUT7 CM_n_net_0.IN a_27642_n32662# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4023 a_35464_5202# a_27682_10411# PRbiased_net_9.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4024 a_29618_n4841# a_27682_n7939# PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4025 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4026 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4027 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4028 PRbiased_net_8.IBN a_47184_10411# a_53562_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4029 PRbiased_net_3.VDD a_47184_n7939# a_47714_n4841# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4030 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4031 a_107014_n10824# PRbiased_net_0.IBN a_106442_n6773# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4032 a_60849_n13906# a_58923_n13906# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4033 a_42168_n38044# CM_n_net_0.IN a_43042_n36250# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4034 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4035 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4036 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4037 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4038 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4039 a_86091_10096# PRbiased_net_6.IBN a_88067_2963# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4040 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4041 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4042 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4043 a_72830_n8314# a_78559_n14221# a_80485_n14221# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4044 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4045 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4046 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4047 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4048 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4049 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4050 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4051 a_29636_n22894# CM_n_net_0.IN a_29076_n21997# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4052 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4053 a_99756_2963# a_97830_2963# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4054 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4055 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4056 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4057 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4058 a_73198_2963# a_66820_10096# a_72676_2963# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4059 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4060 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4061 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4062 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4063 PRbiased_net_2.VDD a_66820_n8254# a_67350_n8254# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4064 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4065 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4066 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4067 FC_top_0.AVDD FC_top_0.IREF a_n11312_n20927# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4068 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4069 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4070 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4071 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4072 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4073 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4074 a_42168_n27379# CM_n_net_0.IN a_43042_n25585# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4075 a_39421_3278# a_39421_3278# a_41347_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4076 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4077 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4078 a_53570_n37186# CM_p_net_0.IN a_52732_n34471# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4079 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4080 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4081 a_n11312_n21934# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4082 PRbiased_net_2.VDD a_66820_n8254# a_67350_n6322# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4083 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4084 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4085 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4086 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4087 a_66992_2903# a_66820_10096# a_73198_6045# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4088 a_86663_2963# a_86263_2903# a_86091_8930# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4089 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4090 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4091 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4092 PRbiased_net_8.IBP a_53194_9185# a_55000_11177# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4093 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4094 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4095 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4096 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4097 a_5821_n12405# a_n11312_n21934# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4098 PRbiased_net_7.VB a_72830_8870# a_74636_8930# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4099 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4100 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4101 a_63560_n20096# CM_p_net_0.IN a_62992_n20096# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4102 a_5821_n12405# a_n11312_n21934# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4103 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4104 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4105 a_34092_9245# a_33692_9185# PRbiased_net_9.VA PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4106 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4107 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4108 a_42168_n33559# CM_n_net_0.IN a_41608_n33559# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4109 a_52164_n39901# CM_p_net_0.IN a_51596_n39901# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4110 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4111 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4112 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4113 a_43042_n39838# CM_n_net_0.IN a_40734_n39838# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4114 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4115 FC_top_0.AVSS a_118181_3278# a_118703_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4116 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4117 a_n540_n22863# a_n10892_n26881# a_n1108_n22863# FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X4118 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4119 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4120 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4121 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4122 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4123 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4124 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4125 a_64128_n34471# CM_p_net_0.IN a_63560_n34471# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4126 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4127 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4128 a_59268_n37186# CM_p_net_0.IN a_58430_n34471# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4129 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4130 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4131 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4132 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4133 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4134 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4135 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4136 a_62154_n25526# CM_p_net_0.IN a_61624_n26431# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4137 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4138 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4139 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4140 a_57294_n25526# CM_p_net_0.IN a_56456_n25526# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4141 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4142 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4143 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4144 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4145 a_50758_n39901# CM_p_net_0.IN a_50228_n39901# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4146 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4147 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4148 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4149 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X4150 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4151 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4152 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4153 a_36776_n39838# CM_n_net_0.IN a_34468_n39838# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4154 a_42168_n22894# CM_n_net_0.IN a_41608_n22894# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4155 a_114224_n11982# a_106442_n6773# PRbiased_net_0.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4156 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4157 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4158 a_93907_8930# a_92101_8870# a_91947_6045# PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4159 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4160 a_92469_n14221# a_86091_n7088# a_91947_n14221# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4161 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4162 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4163 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4164 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4165 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4166 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4167 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4168 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4169 a_108378_9245# a_106442_9245# PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4170 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4171 a_99756_n11139# a_97830_n14221# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4172 a_n1108_n23588# a_n10892_n26881# a_n1676_n23588# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X4173 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4174 FC_top_0.AVDD FC_top_0.IREF a_n11312_n21934# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4175 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4176 PRbiased_net_6.IBN a_86091_10096# a_92469_4887# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4177 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4178 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4179 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4180 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4181 a_118703_3278# a_118181_3278# a_118181_3278# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4182 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4183 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4184 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4185 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4186 PRbiased_net_4.ITP a_27854_n13966# a_39972_n6007# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4187 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4188 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4189 a_49160_5202# PRbiased_net_8.IBN PRbiased_net_8.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4190 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4191 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4192 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4193 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4194 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4195 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4196 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4197 a_40174_n39838# CM_n_net_0.IN a_39652_n39838# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4198 PRbiased_net_7.IBN a_66820_10096# a_73198_4121# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4199 a_31070_n38044# CM_n_net_0.IN a_30510_n38044# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4200 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4201 a_33692_n7999# a_39421_n13906# a_41347_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4202 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4203 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4204 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4205 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4206 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4207 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4208 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4209 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4210 a_80516_10862# PRbiased_net_7.IBP PRbiased_net_7.ITP PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4211 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4212 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4213 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4214 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4215 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4216 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4217 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4218 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4219 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4220 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4221 a_41347_3278# a_39421_3278# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4222 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4223 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4224 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4225 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4226 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4227 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4228 FC_top_0.AVSS a_n11312_n20927# a_n10892_n26881# FC_top_0.AVSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X4229 FC_top_0.AVSS a_72830_8870# a_73230_10862# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4230 a_52732_n38996# CM_p_net_0.IN a_52164_n38996# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4231 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4232 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4233 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4234 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4235 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4236 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4237 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4238 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4239 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4240 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4241 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4242 a_62154_n33566# CM_p_net_0.IN a_61624_n34471# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4243 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4244 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4245 a_57294_n33566# CM_p_net_0.IN a_56456_n33566# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4246 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4247 a_63560_n21001# CM_p_net_0.IN a_62992_n21001# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4248 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4249 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4250 a_27682_9245# a_27854_3218# a_29658_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4251 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4252 a_86263_2903# a_86091_10096# a_92469_2963# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4253 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4254 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4255 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4256 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4257 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4258 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4259 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4260 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4261 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4262 a_28254_n12748# PRbiased_net_4.IBN a_27682_n6773# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4263 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4264 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4265 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4266 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4267 a_108378_n7939# a_106442_n7939# PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4268 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4269 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4270 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4271 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4272 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4273 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4274 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4275 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4276 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4277 a_43602_n35353# CM_n_net_0.IN a_43042_n35353# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4278 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4279 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4280 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4281 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4282 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4283 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4284 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4285 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4286 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4287 a_73230_n7088# a_72830_n8314# PRbiased_net_2.IBP PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4288 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4289 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4290 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4291 a_62154_n24621# CM_p_net_0.IN a_61624_n28241# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4292 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4293 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4294 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4295 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4296 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4297 a_106442_n6773# PRbiased_net_0.IBN a_108418_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4298 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4299 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4300 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4301 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4302 a_n1108_n22863# a_n10892_n26881# a_n1676_n22863# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X4303 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4304 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4305 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4306 a_27682_n6773# a_27682_n7939# a_29618_n7939# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4307 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4308 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4309 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4310 a_n11312_n21934# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4311 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4312 a_118181_3278# a_118181_3278# a_120107_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4313 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4314 a_73230_n5156# a_72830_n8314# PRbiased_net_2.VB PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4315 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4316 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4317 a_28254_4436# PRbiased_net_9.IBN a_27682_10411# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4318 PRbiased_net_5.ITP a_106614_3218# a_118732_9245# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4319 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4320 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4321 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4322 a_47184_9245# a_47184_9245# a_49120_12343# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4323 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4324 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4325 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4326 a_37336_n29173# CM_n_net_0.IN a_36776_n28276# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4327 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4328 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4329 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4330 a_98381_10096# PRbiased_net_6.IBP a_92101_8870# PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4331 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4332 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4333 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4334 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4335 a_53194_n7999# PRbiased_net_3.IBP a_60880_n7939# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4336 a_106972_11177# a_106442_9245# a_106442_9245# PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4337 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4338 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4339 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4340 FC_top_0.AVSS a_118181_3278# a_118703_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4341 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4342 a_66992_n14281# a_66820_n7088# a_73198_n11139# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4343 a_31070_n33559# CM_n_net_0.IN a_30510_n33559# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4344 a_47184_9245# a_47184_9245# a_49120_10411# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4345 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4346 PRbiased_net_3.ITN a_47356_n13966# a_47756_n13906# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4347 PRbiased_net_3.IBN a_47184_n6773# a_53562_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4348 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4349 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4350 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4351 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4352 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4353 a_42168_n33559# CM_n_net_0.IN a_41608_n32662# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4354 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4355 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4356 PRbiased_net_5.ITP PRbiased_net_5.IBP a_118732_12343# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4357 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4358 a_43042_n38941# CM_n_net_0.IN a_42520_n38941# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4359 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4360 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4361 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4362 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4363 a_n13565_n11419# a_n11312_n21934# FC_top_0.VOUT FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4364 PRbiased_net_9.VDD a_27682_9245# a_28212_11177# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4365 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4366 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4367 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4368 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4369 a_n13565_n11419# a_n11312_n21934# FC_top_0.VOUT FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4370 a_86621_10862# a_86091_8930# a_86091_8930# PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4371 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4372 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4373 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4374 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4375 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4376 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4377 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4378 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4379 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4380 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4381 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4382 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4383 a_28254_n10824# PRbiased_net_4.IBN a_27682_n6773# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4384 a_74636_8930# a_72830_8870# a_72676_6045# PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4385 PRbiased_net_5.ITP PRbiased_net_5.IBP a_118732_10411# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4386 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4387 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4388 a_31070_n22894# CM_n_net_0.IN a_30510_n22894# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4389 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4390 a_50758_n24621# CM_p_net_0.IN a_50228_n23716# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4391 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4392 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4393 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4394 a_36776_n38941# CM_n_net_0.IN a_36254_n38941# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4395 a_33908_n27379# CM_n_net_0.IN a_33386_n27379# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4396 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4397 a_47184_10411# PRbiased_net_8.IBN a_49160_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4398 a_118703_5202# a_118181_3278# a_118181_3278# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4399 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4400 PRbiased_net_7.IBN a_66820_10096# a_73198_4887# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4401 a_78559_n14221# a_66992_n14281# a_80516_n7088# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4402 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4403 a_52164_n38091# CM_p_net_0.IN a_51596_n38091# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4404 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4405 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4406 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4407 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4408 a_52732_n39901# CM_p_net_0.IN a_52164_n39901# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4409 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4410 PRbiased_net_6.ITP a_86263_2903# a_98381_10862# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4411 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4412 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4413 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4414 PRbiased_net_0.IBN a_106442_n6773# a_112820_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4415 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4416 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4417 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4418 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4419 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4420 a_47184_n7939# a_47356_n13966# a_49160_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4421 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4422 a_74636_10096# a_72830_8870# FC_top_0.AVSS PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4423 a_59445_6360# a_58923_3278# a_53194_9185# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4424 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4425 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4426 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4427 a_78559_n14221# a_66992_n14281# a_80516_n5156# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4428 a_62154_n32661# CM_p_net_0.IN CM_p_net_0.OUT11 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4429 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4430 PRbiased_net_2.ITP PRbiased_net_2.IBP a_79110_n7088# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4431 a_50758_n38091# CM_p_net_0.IN a_50228_n38091# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4432 a_57294_n32661# CM_p_net_0.IN a_56456_n32661# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4433 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4434 a_40174_n38941# CM_n_net_0.IN a_39652_n39838# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4435 a_57862_n25526# CM_p_net_0.IN a_57294_n25526# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4436 a_43042_n29173# CM_n_net_0.IN a_40734_n29173# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4437 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4438 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4439 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4440 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4441 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4442 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4443 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4444 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4445 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4446 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4447 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4448 a_66820_n8254# a_66992_n14281# a_68796_n13063# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4449 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4450 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4451 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4452 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4453 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4454 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4455 a_66820_10096# a_66820_8930# a_68756_10862# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4456 PRbiased_net_2.ITP PRbiased_net_2.IBP a_79110_n5156# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4457 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4458 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4459 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4460 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4461 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4462 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4463 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4464 a_41347_5202# a_39421_3278# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4465 a_86263_n14281# a_86091_n7088# a_92469_n11139# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4466 a_56456_n25526# CM_p_net_0.IN a_55926_n26431# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4467 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4468 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4469 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4470 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4471 a_36776_n29173# CM_n_net_0.IN a_34468_n29173# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4472 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4473 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4474 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4475 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4476 a_62992_n38996# CM_p_net_0.IN a_62154_n38996# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4477 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4478 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4479 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4480 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4481 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4482 PRbiased_net_6.IBP a_92101_8870# a_93907_10862# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4483 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4484 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4485 a_52164_n31756# CM_p_net_0.IN a_51596_n31756# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4486 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4487 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4488 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4489 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4490 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4491 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4492 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4493 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4494 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4495 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4496 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4497 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4498 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4499 a_40734_n28276# CM_n_net_0.IN a_40174_n28276# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4500 a_112452_n7999# a_118181_n13906# a_120107_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4501 a_55000_9245# a_53194_9185# a_53040_6360# PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4502 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4503 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4504 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4505 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4506 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4507 a_66992_2903# a_66820_10096# a_73198_2963# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4508 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4509 a_106442_9245# a_106614_3218# a_108418_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4510 a_40174_n29173# CM_n_net_0.IN a_39652_n29173# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4511 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4512 a_53594_n6773# a_53194_n7999# PRbiased_net_3.IBP PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4513 a_47756_n11982# a_47356_n13966# a_47184_n7939# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4514 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4515 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4516 a_50758_n31756# CM_p_net_0.IN a_50228_n35376# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4517 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4518 a_106614_n13966# a_106442_n6773# a_112820_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4519 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4520 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4521 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4522 a_67350_n8254# a_66820_n8254# a_66820_n8254# PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4523 a_47184_n7939# a_47356_n13966# a_49160_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4524 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4525 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4526 a_52164_n22811# CM_p_net_0.IN a_51596_n22811# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4527 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4528 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4529 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4530 a_34468_n28276# CM_n_net_0.IN a_33908_n28276# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4531 a_53594_n4841# a_53194_n7999# PRbiased_net_3.VB PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4532 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4533 a_37336_n38044# CM_n_net_0.IN a_36776_n38044# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4534 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4535 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4536 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4537 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4538 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4539 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4540 a_67350_n6322# a_66820_n8254# a_66820_n8254# PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4541 a_28202_n39838# CM_n_net_0.IN a_27642_n39838# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4542 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4543 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4544 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4545 FC_top_0.AVSS a_78559_n14221# a_79081_n11139# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4546 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4547 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4548 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4549 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4550 a_50758_n22811# CM_p_net_0.IN a_50228_n22811# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4551 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4552 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4553 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X4554 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4555 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4556 a_57862_n33566# CM_p_net_0.IN a_57294_n33566# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4557 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4558 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4559 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4560 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4561 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4562 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4563 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4564 a_108418_4436# a_106614_3218# PRbiased_net_5.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4565 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4566 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4567 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4568 a_112298_3278# a_112452_9185# a_112852_9245# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4569 a_120138_12343# a_106614_3218# PRbiased_net_5.ITP PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4570 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4571 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4572 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4573 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4574 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4575 FC_top_0.AVSS a_39421_3278# a_39943_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4576 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4577 a_112852_n7939# a_112452_n7999# PRbiased_net_0.VA PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4578 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4579 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4580 a_64966_n25526# CM_p_net_0.IN a_64128_n25526# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4581 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4582 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4583 PRbiased_net_2.VDD a_66820_n8254# a_67350_n7088# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4584 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4585 a_43042_n24688# CM_n_net_0.IN a_42520_n26482# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4586 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4587 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4588 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4589 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4590 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4591 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4592 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4593 a_108378_n6007# a_106442_n7939# PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4594 a_56456_n33566# CM_p_net_0.IN a_55926_n34471# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4595 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4596 a_120138_10411# a_106614_3218# PRbiased_net_5.ITP PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4597 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4598 a_31070_n33559# CM_n_net_0.IN a_30510_n32662# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4599 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4600 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4601 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4602 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4603 a_118732_9245# a_106614_3218# a_118181_3278# PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4604 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4605 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4606 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4607 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4608 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4609 PRbiased_net_2.VDD a_66820_n8254# a_67350_n5156# PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4610 a_106442_n7939# a_106442_n7939# a_108378_n6773# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4611 a_33908_n37147# CM_n_net_0.IN a_33386_n38044# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4612 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4613 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4614 a_33538_n13906# a_33692_n7999# a_34092_n7939# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4615 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4616 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4617 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4618 a_n11312_n21934# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4619 a_36776_n24688# CM_n_net_0.IN a_36254_n26482# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4620 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4621 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4622 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4623 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4624 a_47184_10411# PRbiased_net_8.IBN a_49160_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4625 a_27682_n6773# a_27682_n7939# a_29618_n6007# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4626 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4627 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4628 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4629 a_47356_3218# a_47184_10411# a_53562_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4630 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4631 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4632 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4633 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4634 a_106442_n7939# a_106442_n7939# a_108378_n4841# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4635 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4636 a_56456_n24621# CM_p_net_0.IN a_55926_n28241# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4637 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4638 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4639 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4640 a_62992_n39901# CM_p_net_0.IN a_62154_n39901# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4641 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4642 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4643 a_60849_n12748# a_58923_n13906# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4644 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4645 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4646 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4647 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4648 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4649 a_78559_n14221# a_78559_n14221# a_80485_n13063# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4650 a_33908_n26482# CM_n_net_0.IN a_33386_n27379# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4651 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4652 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4653 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4654 a_53194_n7999# PRbiased_net_3.IBP a_60880_n6007# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4655 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4656 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4657 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4658 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4659 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4660 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4661 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4662 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4663 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4664 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4665 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4666 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4667 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4668 a_40174_n24688# CM_n_net_0.IN a_39652_n24688# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4669 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4670 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4671 a_n13565_n12405# a_n11312_n21934# a_5821_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4672 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4673 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4674 FC_top_0.AVSS a_97830_n14221# a_98352_n11139# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4675 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4676 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4677 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X4678 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4679 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4680 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4681 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4682 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4683 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4684 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4685 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4686 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4687 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4688 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4689 a_33692_9185# a_39421_3278# a_41347_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4690 a_120107_6360# a_118181_3278# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4691 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4692 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4693 a_86091_8930# a_86091_8930# a_88027_10096# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4694 a_41347_n13906# a_39421_n13906# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4695 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4696 a_37336_n33559# CM_n_net_0.IN a_36776_n33559# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4697 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4698 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4699 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4700 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4701 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4702 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4703 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4704 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4705 a_52732_n38091# CM_p_net_0.IN a_52164_n38091# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4706 a_n1676_n22277# a_n10892_n26881# a_n2206_n22277# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X4707 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4708 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4709 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4710 a_64966_n33566# CM_p_net_0.IN a_64128_n33566# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4711 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4712 a_73230_12028# a_72830_8870# PRbiased_net_7.VB PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4713 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4714 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4715 a_40734_n38941# CM_n_net_0.IN a_40174_n38044# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4716 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4717 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4718 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4719 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4720 PRbiased_net_1.VDD a_86091_n7088# a_93873_n12297# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4721 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4722 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4723 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4724 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X4725 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4726 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4727 a_49120_n6773# a_47184_n7939# PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4728 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4729 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4730 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4731 a_107014_6360# PRbiased_net_5.IBN a_106442_10411# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4732 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4733 PRbiased_net_9.VDD a_27682_9245# a_28212_9245# PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4734 a_41378_n7939# PRbiased_net_4.IBP PRbiased_net_4.ITP PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4735 a_37336_n22894# CM_n_net_0.IN a_36776_n22894# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4736 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4737 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4738 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4739 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4740 a_57862_n32661# CM_p_net_0.IN a_57294_n32661# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4741 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4742 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4743 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4744 a_58430_n25526# CM_p_net_0.IN a_57862_n25526# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4745 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4746 a_91947_n14221# a_92101_n8314# a_92501_n8254# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4747 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4748 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4749 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4750 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4751 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4752 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4753 a_49120_n4841# a_47184_n7939# PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4754 a_60849_n10824# a_58923_n13906# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4755 a_34468_n38941# CM_n_net_0.IN a_33908_n38044# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4756 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4757 a_64966_n24621# CM_p_net_0.IN CM_p_net_0.OUT6 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4758 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4759 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4760 a_92469_n13063# a_86091_n7088# PRbiased_net_1.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4761 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4762 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4763 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4764 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4765 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4766 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4767 a_56456_n32661# CM_p_net_0.IN CM_p_net_0.OUT9 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4768 FC_top_0.AVSS a_92101_n8314# a_92501_n6322# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4769 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4770 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4771 PRbiased_net_9.ITN PRbiased_net_9.IBN a_28254_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4772 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4773 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4774 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4775 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4776 a_63560_n38996# CM_p_net_0.IN a_62992_n38996# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4777 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4778 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4779 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4780 a_39943_4436# a_39421_3278# a_33692_9185# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4781 a_67392_n12297# a_66992_n14281# a_66820_n8254# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4782 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4783 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4784 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4785 a_52732_n31756# CM_p_net_0.IN a_52164_n31756# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4786 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4787 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4788 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4789 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4790 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4791 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X4792 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4793 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4794 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4795 a_33908_n21997# CM_n_net_0.IN a_33386_n22894# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4796 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4797 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4798 a_60880_n7939# PRbiased_net_3.IBP PRbiased_net_3.ITP PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4799 a_92101_n8314# PRbiased_net_1.IBP a_99787_n8254# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4800 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4801 a_28202_n38941# CM_n_net_0.IN a_27642_n38941# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4802 a_43042_n34456# CM_n_net_0.IN a_42520_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4803 a_35464_6360# a_27682_10411# a_27854_3218# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4804 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4805 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4806 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4807 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4808 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4809 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4810 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4811 a_107014_n11982# a_106614_n13966# a_106442_n7939# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4812 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4813 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4814 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4815 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4816 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4817 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4818 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4819 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4820 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4821 a_78559_2963# a_66992_2903# a_80516_12028# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4822 a_92101_n8314# PRbiased_net_1.IBP a_99787_n6322# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4823 a_67350_8930# a_66820_8930# a_66820_8930# PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4824 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4825 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4826 a_35498_n7939# a_33692_n7999# a_33538_n10824# PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4827 a_59474_n7939# a_47356_n13966# a_58923_n13906# PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4828 a_52732_n22811# CM_p_net_0.IN a_52164_n22811# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4829 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4830 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4831 a_n11312_n20927# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X4832 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4833 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4834 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4835 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4836 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4837 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4838 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4839 a_36776_n34456# CM_n_net_0.IN a_36254_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4840 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4841 a_43042_n23791# CM_n_net_0.IN a_42520_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4842 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4843 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4844 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4845 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4846 a_47184_10411# a_47184_9245# a_49120_11177# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4847 PRbiased_net_7.ITP PRbiased_net_7.IBP a_79110_12028# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4848 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4849 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4850 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4851 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4852 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4853 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4854 a_n1676_n21552# a_n10892_n26881# a_n2206_n22277# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X4855 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4856 PRbiased_net_8.IBN a_47184_10411# a_53562_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4857 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4858 a_40734_n34456# CM_n_net_0.IN a_40174_n33559# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4859 a_58430_n33566# CM_p_net_0.IN a_57862_n33566# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4860 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4861 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4862 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4863 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4864 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4865 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4866 a_36776_n23791# CM_n_net_0.IN a_36254_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4867 a_28202_n29173# CM_n_net_0.IN a_27642_n29173# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4868 a_27682_10411# PRbiased_net_9.IBN a_29658_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4869 a_98381_10862# a_86263_2903# a_97830_2963# PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4870 a_40174_n34456# CM_n_net_0.IN a_39652_n35353# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4871 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4872 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4873 a_64966_n33566# CM_p_net_0.IN a_64128_n32661# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4874 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4875 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4876 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4877 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4878 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4879 PRbiased_net_5.ITP a_106614_3218# a_118732_11177# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4880 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4881 a_42168_n39838# CM_n_net_0.IN a_41608_n39838# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4882 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4883 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4884 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4885 a_112852_n6007# a_112452_n7999# PRbiased_net_0.IBP PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4886 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4887 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4888 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4889 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4890 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4891 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4892 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4893 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4894 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4895 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4896 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4897 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4898 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4899 a_34468_n34456# CM_n_net_0.IN a_33908_n33559# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4900 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4901 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4902 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4903 a_40734_n23791# CM_n_net_0.IN a_40174_n22894# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4904 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X4905 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4906 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4907 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4908 FC_top_0.AVSS a_112452_n7999# a_112852_n6773# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4909 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4910 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4911 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4912 a_33692_9185# a_39421_3278# a_41347_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4913 a_40174_n23791# CM_n_net_0.IN a_39652_n24688# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4914 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4915 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4916 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4917 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4918 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4919 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4920 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4921 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4922 a_112452_9185# a_118181_3278# a_120107_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4923 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4924 FC_top_0.AVSS a_n11312_n21934# a_n5714_n27397# FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X4925 a_28254_3278# a_27854_3218# a_27682_9245# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4926 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4927 FC_top_0.AVSS a_33692_n7999# a_34092_n6007# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4928 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4929 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4930 a_112298_n10824# a_112452_n7999# a_112852_n4841# PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4931 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4932 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4933 a_62992_n38091# CM_p_net_0.IN a_62154_n38091# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4934 a_34468_n23791# CM_n_net_0.IN a_33908_n22894# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4935 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4936 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4937 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4938 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4939 a_63560_n39901# CM_p_net_0.IN a_62992_n39901# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4940 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4941 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4942 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4943 a_37336_n33559# CM_n_net_0.IN a_36776_n32662# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4944 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4945 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4946 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4947 a_91947_n11139# a_86091_n7088# a_93873_n14221# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4948 a_99756_n12297# a_97830_n14221# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4949 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4950 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4951 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4952 PRbiased_net_3.ITN PRbiased_net_3.IBN a_47756_n12748# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4953 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4954 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4955 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4956 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4957 a_49160_6360# a_47356_3218# PRbiased_net_8.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4958 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4959 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4960 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4961 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4962 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4963 a_74636_10862# a_72830_8870# FC_top_0.AVSS PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4964 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4965 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4966 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4967 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4968 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4969 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4970 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4971 a_47714_n7939# a_47184_n7939# a_47184_n7939# PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4972 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4973 a_n13565_n12405# a_n11312_n21934# a_5821_n12405# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4974 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4975 a_n13565_n12405# a_n11312_n21934# a_5821_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4976 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4977 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4978 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4979 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4980 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4981 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4982 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4983 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4984 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4985 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4986 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4987 PRbiased_net_7.VDD a_66820_8930# a_67350_12028# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4988 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4989 PRbiased_net_7.VDD a_66820_8930# a_67350_8930# PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4990 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4991 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4992 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4993 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4994 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4995 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4996 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4997 a_67392_n14221# a_66992_n14281# a_66820_n8254# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4998 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4999 PRbiased_net_5.ITN PRbiased_net_5.IBN a_107014_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5000 a_34092_12343# a_33692_9185# PRbiased_net_9.VB PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5001 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5002 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5003 FC_top_0.AVSS a_n11312_n20927# a_n13565_n11419# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5004 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5005 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5006 a_62992_n31756# CM_p_net_0.IN a_62154_n31756# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5007 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5008 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5009 a_51596_n37186# CM_p_net_0.IN a_50758_n37186# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5010 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5011 a_28202_n26482# CM_n_net_0.IN a_27642_n24688# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5012 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5013 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5014 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5015 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5016 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5017 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5018 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5019 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5020 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5021 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5022 a_58430_n32661# CM_p_net_0.IN a_57862_n32661# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5023 a_54966_4436# a_47184_10411# PRbiased_net_8.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5024 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5025 a_34092_10411# a_33692_9185# PRbiased_net_9.IBP PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5026 a_41378_n6007# PRbiased_net_4.IBP PRbiased_net_4.ITP PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5027 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5028 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5029 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5030 a_67350_n7088# a_66820_n8254# a_66820_n7088# PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5031 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5032 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5033 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5034 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5035 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5036 a_39421_n13906# a_27854_n13966# a_41378_n6773# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5037 PRbiased_net_3.ITN PRbiased_net_3.IBN a_47756_n10824# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5038 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5039 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5040 a_30510_n36250# CM_n_net_0.IN a_29636_n34456# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5041 a_62992_n22811# CM_p_net_0.IN a_62154_n22811# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5042 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5043 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5044 a_n11312_n21934# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5045 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5046 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5047 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5048 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5049 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5050 a_51596_n28241# CM_p_net_0.IN a_50758_n28241# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5051 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5052 a_67350_n5156# a_66820_n8254# a_66820_n7088# PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5053 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5054 FC_top_0.AVSS CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5055 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5056 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5057 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5058 a_47184_10411# a_47184_9245# a_49120_9245# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5059 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5060 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5061 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5062 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5063 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5064 a_39421_n13906# a_27854_n13966# a_41378_n4841# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5065 FC_top_0.AVDD FC_top_0.IREF a_n11312_n21934# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5066 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5067 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5068 a_35902_n29173# CM_n_net_0.IN a_35342_n28276# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5069 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5070 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5071 PRbiased_net_3.VB a_53194_n7999# a_55000_n7939# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5072 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5073 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5074 a_72676_2963# a_66820_10096# a_74602_6045# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5075 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5076 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5077 a_120138_11177# PRbiased_net_5.IBP PRbiased_net_5.ITP PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5078 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5079 a_30510_n25585# CM_n_net_0.IN a_29636_n23791# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5080 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5081 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5082 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5083 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5084 a_27682_10411# PRbiased_net_9.IBN a_29658_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5085 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5086 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5087 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5088 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5089 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5090 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5091 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5092 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5093 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5094 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5095 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5096 a_60880_n6007# PRbiased_net_3.IBP PRbiased_net_3.ITP PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5097 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5098 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5099 a_106442_10411# PRbiased_net_5.IBN a_108418_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5100 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5101 CM_n_net_0.OUT11 CM_n_net_0.IN a_40174_n32662# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5102 a_n1676_n23588# a_n10892_n26881# a_n2206_n23588# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X5103 a_29636_n29173# CM_n_net_0.IN a_29076_n28276# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5104 a_n13565_2223# FC_top_0.VP a_n13565_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5105 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5106 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5107 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5108 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5109 FC_top_0.AVSS a_118181_3278# a_118703_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5110 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5111 a_31070_n39838# CM_n_net_0.IN a_30510_n39838# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5112 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5113 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5114 PRbiased_net_2.IBN a_66820_n7088# a_73198_n12297# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5115 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5116 a_118181_3278# a_106614_3218# a_120138_12343# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5117 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5118 a_27642_n36250# CM_n_net_0.IN CM_n_net_0.OUT8 FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5119 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5120 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5121 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5122 a_35498_n6007# a_33692_n7999# FC_top_0.AVSS PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5123 a_42168_n39838# CM_n_net_0.IN a_41608_n38941# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5124 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5125 a_59474_n6007# a_47356_n13966# a_58923_n13906# PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5126 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5127 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5128 a_74602_n11139# a_66820_n7088# a_66992_n14281# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5129 a_51596_n21906# CM_p_net_0.IN a_50758_n21906# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5130 a_74602_6045# a_66820_10096# a_66992_2903# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5131 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5132 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5133 CM_n_net_0.OUT9 CM_n_net_0.IN a_33908_n32662# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5134 a_28254_5202# a_27854_3218# a_27682_9245# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5135 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5136 a_112452_9185# a_118181_3278# a_120107_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5137 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5138 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5139 a_118181_3278# a_106614_3218# a_120138_10411# PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5140 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5141 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5142 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5143 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5144 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5145 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5146 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5147 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5148 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5149 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5150 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5151 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5152 a_28254_n11982# a_27854_n13966# a_27682_n7939# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5153 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5154 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5155 a_27642_n25585# CM_n_net_0.IN CM_n_net_0.OUT2 FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5156 a_108418_3278# PRbiased_net_5.IBN PRbiased_net_5.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5157 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5158 a_68756_10096# a_66820_8930# PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5159 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5160 a_99756_n14221# a_97830_n14221# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5161 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5162 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5163 FC_top_0.AVSS a_39421_3278# a_39943_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5164 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5165 a_118703_6360# a_118181_3278# a_112452_9185# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5166 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5167 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5168 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5169 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5170 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5171 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5172 PRbiased_net_7.VDD a_66820_10096# a_74602_4121# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5173 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5174 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5175 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5176 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5177 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5178 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5179 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5180 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5181 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5182 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5183 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5184 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5185 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5186 a_42168_n29173# CM_n_net_0.IN a_41608_n29173# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5187 a_114258_9245# a_112452_9185# a_112298_6360# PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5188 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5189 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5190 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5191 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5192 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5193 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5194 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5195 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5196 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5197 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5198 a_86091_10096# a_86091_8930# a_88027_10862# PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5199 a_n5714_n26774# a_n11312_n21934# a_n6236_n27397# FC_top_0.AVSS nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X5200 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5201 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5202 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5203 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5204 a_63560_n38091# CM_p_net_0.IN a_62992_n38091# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5205 a_28202_n34456# CM_n_net_0.IN a_27642_n34456# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5206 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5207 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5208 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5209 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5210 a_41347_6360# a_39421_3278# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5211 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5212 PRbiased_net_1.IBN a_86091_n7088# a_92469_n12297# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5213 a_74602_4121# a_66820_10096# PRbiased_net_7.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5214 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5215 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5216 FC_top_0.AVSS a_92101_n8314# a_92501_n7088# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5217 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5218 a_n1676_n22863# a_n10892_n26881# a_n2206_n23588# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X5219 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5220 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5221 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5222 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5223 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5224 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5225 a_53040_6360# a_53194_9185# a_53594_12343# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5226 a_28202_n23791# CM_n_net_0.IN a_27642_n23791# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5227 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5228 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5229 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5230 a_91947_n11139# a_92101_n8314# a_92501_n5156# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5231 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5232 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5233 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5234 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5235 a_47714_n6007# a_47184_n7939# a_47184_n7939# PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5236 a_53570_n37186# CM_p_net_0.IN a_52732_n37186# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5237 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5238 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5239 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5240 a_41347_n12748# a_39421_n13906# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5241 a_43602_n27379# CM_n_net_0.IN a_43042_n27379# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5242 FC_top_0.AVSS a_53194_9185# a_53594_10411# PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5243 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5244 a_35902_n38044# CM_n_net_0.IN a_35342_n38044# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5245 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5246 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5247 PRbiased_net_0.IBN a_106442_n6773# a_112820_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5248 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5249 a_47184_n6773# PRbiased_net_3.IBN a_49160_n11982# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5250 a_30510_n35353# CM_n_net_0.IN a_29988_n37147# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5251 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5252 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5253 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5254 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5255 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5256 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5257 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5258 a_63560_n31756# CM_p_net_0.IN a_62992_n31756# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5259 a_97830_n14221# a_86263_n14281# a_99787_n7088# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5260 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5261 a_106972_n7939# a_106442_n7939# a_106442_n7939# PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5262 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5263 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5264 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5265 a_64128_n37186# CM_p_net_0.IN a_63560_n37186# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5266 a_29636_n38044# CM_n_net_0.IN a_29076_n38044# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5267 FC_top_0.AVSS a_78559_n14221# a_79081_n12297# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5268 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5269 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5270 CM_p_net_0.VDD CM_p_net_0.IN a_52732_n28241# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5271 a_59268_n37186# CM_p_net_0.IN a_58430_n37186# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5272 a_106442_10411# PRbiased_net_5.IBN a_108418_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5273 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5274 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5275 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5276 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5277 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5278 a_97830_n14221# a_86263_n14281# a_99787_n5156# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5279 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5280 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5281 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5282 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5283 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5284 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5285 a_n11312_n20927# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5286 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5287 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5288 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5289 a_66992_n14281# a_66820_n7088# a_73198_n14221# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5290 a_63560_n22811# CM_p_net_0.IN a_62992_n22811# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5291 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5292 a_92469_6045# a_86091_10096# a_91947_6045# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5293 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5294 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5295 PRbiased_net_4.VDD a_27682_n7939# a_28212_n7939# PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5296 CM_n_net_0.IN CM_n_net_0.IN FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5297 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5298 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5299 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5300 PRbiased_net_9.ITN a_27854_3218# a_28254_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5301 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5302 a_64128_n28241# CM_p_net_0.IN a_63560_n28241# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5303 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5304 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X5305 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5306 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5307 a_31070_n39838# CM_n_net_0.IN a_30510_n38941# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5308 CM_p_net_0.VDD CM_p_net_0.IN a_58430_n28241# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5309 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5310 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5311 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5312 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5313 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5314 a_27642_n35353# CM_n_net_0.IN a_27120_n35353# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5315 FC_top_0.AVDD FC_top_0.IREF a_n11312_n21934# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5316 a_39943_3278# a_39421_3278# a_39421_3278# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5317 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5318 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5319 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5320 a_n13565_n11419# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5321 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5322 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5323 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5324 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5325 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5326 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5327 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5328 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5329 PRbiased_net_3.IBP a_53194_n7999# a_55000_n6007# PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5330 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5331 a_108418_5202# PRbiased_net_5.IBN PRbiased_net_5.ITN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5332 a_41347_n10824# a_39421_n13906# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5333 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5334 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5335 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5336 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5337 PRbiased_net_7.VDD a_66820_10096# a_74602_4887# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5338 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5339 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5340 a_47714_9245# a_47184_9245# a_47184_9245# PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5341 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5342 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5343 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5344 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5345 FC_top_0.AVSS a_n11312_n20927# a_n13565_n12405# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5346 FC_top_0.AVSS a_39421_3278# a_39943_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5347 a_47184_9245# a_47356_3218# a_49160_6360# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5348 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5349 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5350 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5351 a_53570_n21906# CM_p_net_0.IN a_52732_n21906# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5352 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5353 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5354 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5355 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5356 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5357 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5358 a_86091_n8254# a_86263_n14281# a_88067_n11139# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5359 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5360 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5361 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5362 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5363 a_n13565_n11419# a_n11312_n21934# FC_top_0.VOUT FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5364 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5365 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5366 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5367 FC_top_0.VOUT a_n10892_n26881# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5368 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5369 a_80516_8930# PRbiased_net_7.IBP PRbiased_net_7.ITP PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5370 a_n13565_n11419# FC_top_0.VN a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5371 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5372 a_51596_n20096# CM_p_net_0.IN a_50758_n20096# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5373 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5374 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5375 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5376 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5377 a_35902_n33559# CM_n_net_0.IN a_35342_n33559# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5378 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5379 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5380 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5381 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5382 FC_top_0.AVSS a_97830_n14221# a_98352_n12297# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5383 a_31070_n29173# CM_n_net_0.IN a_30510_n29173# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5384 a_n13565_n12405# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5385 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5386 a_64128_n21906# CM_p_net_0.IN a_63560_n21906# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5387 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5388 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5389 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5390 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5391 a_74602_4887# a_66820_10096# PRbiased_net_7.IBN FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5392 a_93907_n8254# a_92101_n8314# a_91947_n11139# PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5393 a_53570_n36281# CM_p_net_0.IN CM_p_net_0.OUT8 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5394 a_59268_n21906# CM_p_net_0.IN a_58430_n21906# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5395 a_67350_12028# a_66820_8930# a_66820_10096# PRbiased_net_7.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5396 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5397 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5398 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5399 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5400 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5401 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5402 a_92469_4121# a_86091_10096# PRbiased_net_6.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5403 a_37336_n39838# CM_n_net_0.IN a_36776_n39838# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5404 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5405 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5406 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5407 a_86263_n14281# a_86091_n7088# a_92469_n14221# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5408 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5409 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5410 a_35464_n13906# a_27682_n6773# a_27854_n13966# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5411 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5412 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5413 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5414 a_29636_n33559# CM_n_net_0.IN a_29076_n33559# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5415 a_5821_3209# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5416 PRbiased_net_8.VDD a_47184_10411# a_54966_4436# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5417 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5418 a_93907_n6322# a_92101_n8314# FC_top_0.AVSS PRbiased_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5419 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5420 a_97830_n14221# a_97830_n14221# a_99756_n11139# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5421 a_35902_n22894# CM_n_net_0.IN a_35342_n22894# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5422 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5423 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5424 a_n13565_2223# FC_top_0.VN a_n13565_n11419# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5425 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5426 PRbiased_net_1.VDD a_86091_n8254# a_86621_n8254# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5427 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5428 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5429 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5430 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5431 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5432 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5433 FC_top_0.AVDD FC_top_0.IREF a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5434 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5435 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5436 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5437 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5438 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5439 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5440 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5441 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5442 a_43602_n38044# CM_n_net_0.IN a_43042_n37147# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5443 a_59268_n36281# CM_p_net_0.IN CM_p_net_0.OUT10 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5444 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5445 a_72676_6045# a_66820_10096# a_74602_2963# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5446 a_62154_n27336# CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5447 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5448 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5449 PRbiased_net_1.VDD a_86091_n8254# a_86621_n6322# PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5450 a_57294_n27336# CM_p_net_0.IN a_56456_n27336# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5451 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5452 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5453 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5454 a_29636_n22894# CM_n_net_0.IN a_29076_n22894# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5455 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5456 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5457 a_5821_2223# a_n10892_n26881# a_5821_n12405# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5458 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5459 a_60849_n11982# a_58923_n13906# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5460 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5461 a_34092_11177# a_33692_9185# PRbiased_net_9.IBP PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5462 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5463 a_53562_4436# a_47184_10411# PRbiased_net_8.VDD FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5464 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5465 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5466 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5467 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5468 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5469 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5470 a_5821_2223# a_5821_n12405# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5471 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5472 a_43602_n27379# CM_n_net_0.IN a_43042_n26482# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5473 a_39972_n6773# PRbiased_net_4.IBP a_33692_n7999# PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5474 PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD PRbiased_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5475 PRbiased_net_1.VDD a_86091_n7088# a_93873_n13063# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5476 FC_top_0.AVDD a_5821_n12405# a_5821_3209# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5477 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5478 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5479 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5480 a_59445_n13906# a_58923_n13906# a_58923_n13906# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5481 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5482 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5483 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5484 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5485 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5486 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5487 FC_top_0.AVSS a_78559_n14221# a_79081_n14221# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5488 a_74602_2963# a_66820_10096# a_66992_2903# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5489 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5490 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5491 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5492 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5493 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5494 a_39972_n4841# PRbiased_net_4.IBP a_33692_n7999# PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5495 a_n5714_n26221# a_n11312_n21934# a_n11312_n21934# FC_top_0.AVSS nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X5496 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5497 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5498 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5499 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5500 PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD PRbiased_net_3.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5501 a_n10892_n26881# a_n11312_n20927# FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X5502 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5503 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5504 a_5821_n12405# a_n10892_n26881# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5505 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5506 a_42168_n34456# CM_n_net_0.IN a_41608_n34456# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5507 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5508 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5509 FC_top_0.AVDD a_5821_n12405# a_5821_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5510 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5511 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5512 a_n11312_n21934# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5513 PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD PRbiased_net_5.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5514 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5515 PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD PRbiased_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5516 a_n13565_n12405# FC_top_0.VP a_n13565_2223# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5517 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5518 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5519 a_35342_n27379# CM_n_net_0.IN a_34820_n28276# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5520 PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD PRbiased_net_4.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5521 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5522 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5523 PRbiased_net_9.ITN a_27854_3218# a_28254_5202# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5524 a_31070_n24688# CM_n_net_0.IN a_30510_n24688# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5525 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5526 PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD PRbiased_net_7.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5527 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5528 a_51596_n21001# CM_p_net_0.IN a_50758_n21001# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5529 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5530 PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD PRbiased_net_2.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5531 PRbiased_net_5.ITN a_106614_3218# a_107014_3278# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5532 a_67392_n13063# PRbiased_net_2.IBN a_66820_n7088# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5533 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5534 FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5535 a_n13565_2223# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5536 a_39943_5202# a_39421_3278# a_39421_3278# FC_top_0.AVSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5537 a_42168_n23791# CM_n_net_0.IN a_41608_n23791# FC_top_0.AVSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5538 PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD PRbiased_net_9.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5539 PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD PRbiased_net_8.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5540 a_5821_3209# a_n10892_n26881# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5541 PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD PRbiased_net_6.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
.ends

