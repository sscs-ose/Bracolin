* Extracted by KLayout with GF180MCU LVS runset on : 23/03/2024 07:14

.SUBCKT SAR_Asynchornous_Logic
M$1 VDDD \$45 \$14 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$2 VDDD \$44 \$73 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$3 VDDD \$51 \$44 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$4 \$10 \$73 \$3 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$5 \$108 Set \$10 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$6 VDDD \$45 \$108 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$7 \$109 \$3 \$45 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$8 VDDD \$46 \$109 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$9 \$11 \$44 \$3 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$10 \$12 \$44 \$9 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$11 \$110 \$46 \$12 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$12 VDDD \$11 \$110 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$13 \$111 \$9 \$11 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$14 VDDD Set \$111 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$15 \$15 \$73 \$9 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$16 \$16 \$47 \$15 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$17 \$47 CLK VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$18 VSSD \$47 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$19 \$177 \$215 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$20 \$178 \$177 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$21 \$172 \$178 \$171 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$22 \$280 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$23 \$173 \$172 \$280 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$24 \$281 \$173 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$25 \$174 \$46 \$281 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$26 \$172 \$177 \$174 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$27 \$176 \$177 \$173 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$28 \$282 \$46 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$29 \$15 \$176 \$282 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$30 \$283 \$15 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$31 \$175 Set \$283 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$32 \$176 \$178 \$175 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$33 \$179 \$15 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$34 \$15 VSSD VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$35 \$16 \$241 \$15 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$36 \$13 \$15 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$37 \$180 VSSD \$13 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$38 VSSD \$15 \$13 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$39 \$15 \$47 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$40 \$16 VSSD \$15 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$41 \$10 \$44 \$3 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$42 \$10 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$43 VSSD \$45 \$10 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$44 \$45 \$3 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$45 VSSD \$46 \$45 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$46 \$11 \$73 \$3 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$47 \$12 \$73 \$9 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$48 \$12 \$46 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$49 VSSD \$11 \$12 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$50 \$11 \$9 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$51 VSSD Set \$11 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$52 \$15 \$44 \$9 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$53 VSSD \$45 \$14 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$54 \$172 \$177 \$171 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$55 \$173 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$56 VSSD \$172 \$173 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$57 \$174 \$173 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$58 VSSD \$46 \$174 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$59 \$172 \$178 \$174 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$60 \$176 \$178 \$173 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$61 \$15 \$46 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$62 VSSD \$176 \$15 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$63 \$175 \$15 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$64 VSSD Set \$175 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$65 \$176 \$177 \$175 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$66 VSSD \$44 \$73 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$67 VSSD \$51 \$44 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$68 \$47 CLK VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$69 VSSD \$47 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$70 \$177 \$215 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$71 \$178 \$177 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$72 \$179 \$15 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$73 \$16 VSSD \$15 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$74 \$180 \$47 \$13 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
.ENDS SAR_Asynchornous_Logic
