* Extracted by KLayout with GF180MCU LVS runset on : 02/04/2024 15:15

.SUBCKT Filter_TOP VCM IN_POS VDD VSS OUT IBPOUT IBNOUT I1N I1U IN_NEG
M$1 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$4 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$5 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$6 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$7 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$8 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$9 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$10 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$11 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$12 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$13 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$14 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$15 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$16 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$17 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$18 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$19 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$20 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$21 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$22 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$23 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$24 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$25 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$26 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$27 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$28 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$29 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$30 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$31 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$32 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$33 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$34 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$35 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$36 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$37 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$38 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$39 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$40 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$41 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$42 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$43 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$44 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$45 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$46 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$47 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$48 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$49 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$50 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$51 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$52 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$53 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$54 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$55 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$56 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$57 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$58 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$59 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$60 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$61 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$62 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$63 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$64 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$65 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$66 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$67 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$68 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$69 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$70 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$71 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$72 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$73 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$74 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$75 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$76 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$77 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$78 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$79 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$80 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$81 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$82 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$83 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$84 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$85 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$86 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$87 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$88 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$89 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$90 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$91 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$92 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$93 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$94 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$95 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$96 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$97 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$98 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$99 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$100 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$101 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$102 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$103 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$104 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$105 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$106 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$107 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$108 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$109 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$110 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$111 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$112 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$113 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$114 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$115 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$116 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$117 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$118 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$119 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$120 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$121 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$122 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$123 \$145 \$180 \$925 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$124 VDD \$180 \$145 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$125 \$146 \$180 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$126 \$180 \$180 \$146 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$127 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$128 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$129 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$130 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$131 \$147 \$34 \$10 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$132 \$148 \$34 \$147 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$133 \$149 \$34 \$125 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$134 \$6 \$34 \$149 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$135 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$136 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$137 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$138 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$139 \$150 \$181 \$34 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$140 \$39 \$181 \$150 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$141 \$151 \$266 \$39 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$142 \$265 \$266 \$151 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$143 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$144 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$145 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$146 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$147 \$152 \$182 \$927 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$148 VDD \$182 \$152 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$149 \$153 \$182 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$150 \$182 \$182 \$153 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$151 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$152 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$153 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$154 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$155 \$154 \$35 \$11 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$156 \$155 \$35 \$154 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$157 \$156 \$35 \$126 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$158 \$10 \$35 \$156 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$159 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$160 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$161 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$162 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$163 \$157 \$183 \$35 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$164 \$40 \$183 \$157 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$165 \$158 \$268 \$40 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$166 \$267 \$268 \$158 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$167 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$168 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$169 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$170 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$171 \$159 \$184 \$929 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$172 VDD \$184 \$159 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$173 \$160 \$184 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$174 \$184 \$184 \$160 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$175 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$176 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$177 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$178 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$179 \$161 \$36 \$12 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$180 \$162 \$36 \$161 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$181 \$163 \$36 \$127 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$182 \$11 \$36 \$163 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$183 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$184 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$185 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$186 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$187 \$164 \$185 \$36 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$188 \$41 \$185 \$164 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$189 \$165 \$270 \$41 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$190 \$269 \$270 \$165 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$191 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$192 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$193 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$194 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$195 \$166 \$186 \$931 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$196 VDD \$186 \$166 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$197 \$167 \$186 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$198 \$186 \$186 \$167 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$199 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$200 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$201 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$202 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$203 \$168 \$37 \$13 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$204 \$169 \$37 \$168 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$205 \$170 \$37 \$128 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$206 \$12 \$37 \$170 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$207 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$208 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$209 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$210 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$211 \$171 \$187 \$37 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$212 \$42 \$187 \$171 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$213 \$172 \$272 \$42 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$214 \$271 \$272 \$172 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$215 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$216 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$217 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$218 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$219 \$173 \$188 \$933 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$220 VDD \$188 \$173 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$221 \$174 \$188 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$222 \$188 \$188 \$174 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$223 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$224 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$225 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$226 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$227 \$175 \$38 VCM VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$228 \$176 \$38 \$175 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$229 \$177 \$38 \$129 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$230 \$13 \$38 \$177 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$231 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$232 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$233 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$234 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$235 \$178 \$189 \$38 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$236 \$43 \$189 \$178 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$237 \$179 \$274 \$43 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$238 \$273 \$274 \$179 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$239 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$240 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$241 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$242 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$243 \$330 \$180 \$180 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$244 VDD \$180 \$330 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$245 \$331 \$180 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$246 \$925 \$180 \$331 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$247 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$248 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$249 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$250 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$251 \$332 \$34 \$181 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$252 VSS \$34 \$332 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$253 \$333 \$34 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$254 \$181 \$34 \$333 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$255 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$256 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$257 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$258 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$259 \$334 \$266 \$265 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$260 \$39 \$266 \$334 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$261 \$335 \$181 \$39 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$262 \$34 \$181 \$335 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$263 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$264 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$265 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$266 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$267 \$336 \$182 \$182 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$268 VDD \$182 \$336 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$269 \$337 \$182 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$270 \$927 \$182 \$337 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$271 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$272 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$273 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$274 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$275 \$338 \$35 \$183 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$276 VSS \$35 \$338 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$277 \$339 \$35 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$278 \$183 \$35 \$339 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$279 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$280 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$281 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$282 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$283 \$340 \$268 \$267 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$284 \$40 \$268 \$340 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$285 \$341 \$183 \$40 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$286 \$35 \$183 \$341 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$287 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$288 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$289 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$290 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$291 \$342 \$184 \$184 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$292 VDD \$184 \$342 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$293 \$343 \$184 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$294 \$929 \$184 \$343 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$295 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$296 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$297 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$298 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$299 \$344 \$36 \$185 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$300 VSS \$36 \$344 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$301 \$345 \$36 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$302 \$185 \$36 \$345 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$303 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$304 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$305 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$306 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$307 \$346 \$270 \$269 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$308 \$41 \$270 \$346 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$309 \$347 \$185 \$41 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$310 \$36 \$185 \$347 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$311 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$312 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$313 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$314 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$315 \$348 \$186 \$186 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$316 VDD \$186 \$348 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$317 \$349 \$186 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$318 \$931 \$186 \$349 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$319 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$320 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$321 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$322 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$323 \$350 \$37 \$187 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$324 VSS \$37 \$350 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$325 \$351 \$37 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$326 \$187 \$37 \$351 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$327 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$328 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$329 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$330 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$331 \$352 \$272 \$271 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$332 \$42 \$272 \$352 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$333 \$353 \$187 \$42 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$334 \$37 \$187 \$353 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$335 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$336 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$337 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$338 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$339 \$354 \$188 \$188 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$340 VDD \$188 \$354 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$341 \$355 \$188 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$342 \$933 \$188 \$355 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$343 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$344 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$345 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$346 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$347 \$356 \$38 \$189 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$348 VSS \$38 \$356 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$349 \$357 \$38 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$350 \$189 \$38 \$357 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$351 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$352 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$353 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$354 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$355 \$358 \$274 \$273 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$356 \$43 \$274 \$358 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$357 \$359 \$189 \$43 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$358 \$38 \$189 \$359 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$359 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$360 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$361 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$362 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$363 \$450 \$180 \$925 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$364 VDD \$180 \$450 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$365 \$451 \$180 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$366 \$180 \$180 \$451 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$367 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$368 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$369 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$370 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$371 \$452 \$34 \$181 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$372 VSS \$34 \$452 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$373 \$453 \$34 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$374 \$181 \$34 \$453 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$375 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$376 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$377 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$378 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$379 \$454 \$181 \$34 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$380 \$39 \$181 \$454 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$381 \$455 \$266 \$39 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$382 \$265 \$266 \$455 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$383 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$384 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$385 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$386 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$387 \$456 \$182 \$927 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$388 VDD \$182 \$456 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$389 \$457 \$182 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$390 \$182 \$182 \$457 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$391 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$392 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$393 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$394 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$395 \$458 \$35 \$183 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$396 VSS \$35 \$458 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$397 \$459 \$35 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$398 \$183 \$35 \$459 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$399 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$400 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$401 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$402 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$403 \$460 \$183 \$35 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$404 \$40 \$183 \$460 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$405 \$461 \$268 \$40 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$406 \$267 \$268 \$461 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$407 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$408 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$409 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$410 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$411 \$462 \$184 \$929 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$412 VDD \$184 \$462 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$413 \$463 \$184 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$414 \$184 \$184 \$463 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$415 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$416 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$417 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$418 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$419 \$464 \$36 \$185 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$420 VSS \$36 \$464 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$421 \$465 \$36 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$422 \$185 \$36 \$465 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$423 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$424 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$425 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$426 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$427 \$466 \$185 \$36 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$428 \$41 \$185 \$466 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$429 \$467 \$270 \$41 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$430 \$269 \$270 \$467 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$431 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$432 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$433 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$434 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$435 \$468 \$186 \$931 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$436 VDD \$186 \$468 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$437 \$469 \$186 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$438 \$186 \$186 \$469 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$439 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$440 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$441 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$442 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$443 \$470 \$37 \$187 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$444 VSS \$37 \$470 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$445 \$471 \$37 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$446 \$187 \$37 \$471 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$447 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$448 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$449 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$450 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$451 \$472 \$187 \$37 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$452 \$42 \$187 \$472 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$453 \$473 \$272 \$42 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$454 \$271 \$272 \$473 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$455 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$456 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$457 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$458 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$459 \$474 \$188 \$933 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$460 VDD \$188 \$474 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$461 \$475 \$188 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$462 \$188 \$188 \$475 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$463 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$464 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$465 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$466 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$467 \$476 \$38 \$189 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$468 VSS \$38 \$476 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$469 \$477 \$38 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$470 \$189 \$38 \$477 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$471 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$472 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$473 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$474 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$475 \$478 \$189 \$38 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$476 \$43 \$189 \$478 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$477 \$479 \$274 \$43 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$478 \$273 \$274 \$479 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$479 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$480 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$481 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$482 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$483 \$595 \$180 \$180 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$484 VDD \$180 \$595 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$485 \$596 \$180 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$486 \$925 \$180 \$596 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$487 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$488 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$489 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$490 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$491 \$597 \$34 \$6 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$492 \$125 \$34 \$597 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$493 \$598 \$34 \$148 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$494 \$10 \$34 \$598 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$495 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$496 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$497 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$498 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$499 \$599 \$266 \$265 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$500 \$39 \$266 \$599 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$501 \$600 \$181 \$39 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$502 \$34 \$181 \$600 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$503 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$504 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$505 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$506 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$507 \$601 \$182 \$182 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$508 VDD \$182 \$601 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$509 \$602 \$182 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$510 \$927 \$182 \$602 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$511 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$512 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$513 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$514 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$515 \$603 \$35 \$10 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$516 \$126 \$35 \$603 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$517 \$604 \$35 \$155 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$518 \$11 \$35 \$604 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$519 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$520 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$521 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$522 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$523 \$605 \$268 \$267 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$524 \$40 \$268 \$605 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$525 \$606 \$183 \$40 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$526 \$35 \$183 \$606 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$527 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$528 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$529 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$530 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$531 \$607 \$184 \$184 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$532 VDD \$184 \$607 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$533 \$608 \$184 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$534 \$929 \$184 \$608 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$535 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$536 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$537 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$538 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$539 \$609 \$36 \$11 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$540 \$127 \$36 \$609 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$541 \$610 \$36 \$162 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$542 \$12 \$36 \$610 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$543 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$544 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$545 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$546 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$547 \$611 \$270 \$269 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$548 \$41 \$270 \$611 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$549 \$612 \$185 \$41 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$550 \$36 \$185 \$612 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$551 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$552 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$553 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$554 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$555 \$613 \$186 \$186 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$556 VDD \$186 \$613 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$557 \$614 \$186 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$558 \$931 \$186 \$614 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$559 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$560 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$561 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$562 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$563 \$615 \$37 \$12 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$564 \$128 \$37 \$615 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$565 \$616 \$37 \$169 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$566 \$13 \$37 \$616 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$567 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$568 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$569 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$570 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$571 \$617 \$272 \$271 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$572 \$42 \$272 \$617 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$573 \$618 \$187 \$42 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$574 \$37 \$187 \$618 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$575 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$576 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$577 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$578 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$579 \$619 \$188 \$188 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$580 VDD \$188 \$619 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$581 \$620 \$188 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$582 \$933 \$188 \$620 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$583 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$584 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$585 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$586 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$587 \$621 \$38 \$13 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$588 \$129 \$38 \$621 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$589 \$622 \$38 \$176 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$590 VCM \$38 \$622 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$591 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$592 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$593 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$594 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$595 \$623 \$274 \$273 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$596 \$43 \$274 \$623 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$597 \$624 \$189 \$43 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$598 \$38 \$189 \$624 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$599 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$600 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$601 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$602 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$603 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$604 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$605 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$606 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$607 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$608 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$609 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$610 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$611 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$612 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$613 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$614 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$615 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$616 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$617 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$618 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$619 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$620 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$621 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$622 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$623 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$624 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$625 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$626 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$627 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$628 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$629 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$630 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$631 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$632 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$633 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$634 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$635 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$636 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$637 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$638 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$639 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$640 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$641 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$642 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$643 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$644 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$645 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$646 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$647 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$648 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$649 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$650 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$651 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$652 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$653 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$654 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$655 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$656 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$657 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$658 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$659 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$660 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$661 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$662 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$663 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$664 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$665 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$666 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$667 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$668 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$669 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$670 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$671 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$672 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$673 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$674 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$675 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$676 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$677 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$678 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$679 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$680 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$681 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$682 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$683 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$684 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$685 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$686 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$687 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$688 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$689 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$690 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$691 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$692 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$693 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$694 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$695 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$696 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$697 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$698 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$699 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$700 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$701 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$702 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$703 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$704 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$705 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$706 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$707 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$708 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$709 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$710 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$711 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$712 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$713 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$714 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$715 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$716 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$717 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$718 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$719 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$720 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$721 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$722 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$723 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$724 \$1592 \$1581 \$1591 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$725 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$726 \$1679 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$727 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$728 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$729 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$730 \$1593 \$1581 \$1592 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$731 \$1594 \$1581 \$1593 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$732 \$1595 \$1581 \$1594 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$733 \$1680 \$1581 \$1679 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$734 \$1681 \$1581 \$1680 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$735 \$1682 \$1581 \$1681 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$736 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$737 VDD \$1581 \$1595 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$738 \$1683 \$1581 \$1682 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$739 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$740 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$741 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$742 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$743 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$744 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$745 \$1684 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$746 \$1597 \$1581 \$1596 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$747 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$748 \$1598 \$1581 \$1597 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$749 \$1599 \$1581 \$1598 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$750 \$1600 \$1581 \$1599 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$751 \$1685 \$1581 \$1684 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$752 \$1686 \$1581 \$1685 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$753 \$1687 \$1581 \$1686 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$754 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$755 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$756 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$757 VDD \$1581 \$1600 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$758 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$759 \$1688 \$1581 \$1687 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$760 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$761 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$762 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$763 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$764 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$765 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$766 \$1689 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$767 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$768 \$1602 \$1581 \$1601 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$769 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$770 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$771 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$772 \$1603 \$1581 \$1602 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$773 \$1604 \$1581 \$1603 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$774 \$1605 \$1581 \$1604 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$775 \$1690 \$1581 \$1689 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$776 \$1691 \$1581 \$1690 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$777 \$1692 \$1581 \$1691 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$778 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$779 VDD \$1581 \$1605 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$780 \$1693 \$1581 \$1692 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$781 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$782 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$783 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$784 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$785 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$786 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$787 \$1694 \$1582 \$181 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$788 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$789 \$1607 \$1582 \$1606 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$790 \$1695 \$1582 \$1694 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$791 \$1696 \$1582 \$1695 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$792 \$1697 \$1582 \$1696 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$793 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$794 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$795 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$796 \$1608 \$1582 \$1607 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$797 \$1609 \$1582 \$1608 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$798 \$1610 \$1582 \$1609 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$799 \$1611 \$1582 \$1610 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$800 \$1698 \$1582 \$1697 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$801 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$802 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$803 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$804 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$805 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$806 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$807 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$808 \$1699 \$1582 \$183 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$809 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$810 \$1613 \$1582 \$1612 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$811 \$1614 \$1582 \$1613 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$812 \$1615 \$1582 \$1614 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$813 \$1616 \$1582 \$1615 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$814 \$1700 \$1582 \$1699 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$815 \$1701 \$1582 \$1700 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$816 \$1702 \$1582 \$1701 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$817 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$818 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$819 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$820 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$821 \$1617 \$1582 \$1616 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$822 \$1703 \$1582 \$1702 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$823 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$824 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$825 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$826 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$827 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$828 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$829 \$1619 \$1582 \$1618 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$830 \$1704 \$1582 \$185 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$831 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$832 \$1705 \$1582 \$1704 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$833 \$1706 \$1582 \$1705 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$834 \$1707 \$1582 \$1706 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$835 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$836 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$837 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$838 \$1620 \$1582 \$1619 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$839 \$1621 \$1582 \$1620 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$840 \$1622 \$1582 \$1621 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$841 \$1708 \$1582 \$1707 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$842 \$1623 \$1582 \$1622 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$843 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$844 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$845 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$846 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$847 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$848 \$1835 \$1581 \$1834 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$849 \$1836 \$1581 \$1835 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$850 \$1837 \$1581 \$1836 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$851 \$1838 \$1581 \$1837 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$852 \$1683 \$1581 \$1838 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$853 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$854 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$855 \$1840 \$1581 \$1839 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$856 \$1841 \$1581 \$1840 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$857 \$1842 \$1581 \$1841 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$858 \$1843 \$1581 \$1842 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$859 \$1688 \$1581 \$1843 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$860 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$861 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$862 \$1845 \$1581 \$1844 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$863 \$1846 \$1581 \$1845 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$864 \$1847 \$1581 \$1846 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$865 \$1848 \$1581 \$1847 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$866 \$1693 \$1581 \$1848 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$867 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$868 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$869 \$1850 \$1582 \$1849 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$870 \$1851 \$1582 \$1850 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$871 \$1852 \$1582 \$1851 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$872 \$1853 \$1582 \$1852 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$873 \$1698 \$1582 \$1853 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$874 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$875 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$876 \$1855 \$1582 \$1854 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$877 \$1856 \$1582 \$1855 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$878 \$1857 \$1582 \$1856 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$879 \$1858 \$1582 \$1857 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$880 \$1703 \$1582 \$1858 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$881 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$882 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$883 \$1860 \$1582 \$1859 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$884 \$1861 \$1582 \$1860 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$885 \$1862 \$1582 \$1861 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$886 \$1863 \$1582 \$1862 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$887 \$1708 \$1582 \$1863 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$888 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$889 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$890 \$1984 \$1581 \$1834 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$891 \$1985 \$1581 \$1984 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$892 \$1986 \$1581 \$1985 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$893 \$1987 \$1581 \$1986 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$894 \$1988 \$1581 \$1987 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$895 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$896 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$897 \$1989 \$1581 \$1839 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$898 \$1990 \$1581 \$1989 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$899 \$1991 \$1581 \$1990 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$900 \$1992 \$1581 \$1991 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$901 \$1993 \$1581 \$1992 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$902 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$903 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$904 \$1994 \$1581 \$1844 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$905 \$1995 \$1581 \$1994 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$906 \$1996 \$1581 \$1995 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$907 \$1997 \$1581 \$1996 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$908 \$1998 \$1581 \$1997 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$909 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$910 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$911 \$1999 \$1582 \$1849 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$912 \$2000 \$1582 \$1999 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$913 \$2001 \$1582 \$2000 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$914 \$2002 \$1582 \$2001 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$915 \$2003 \$1582 \$2002 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$916 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$917 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$918 \$2004 \$1582 \$1854 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$919 \$2005 \$1582 \$2004 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$920 \$2006 \$1582 \$2005 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$921 \$2007 \$1582 \$2006 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$922 \$2008 \$1582 \$2007 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$923 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$924 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$925 \$2009 \$1582 \$1859 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$926 \$2010 \$1582 \$2009 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$927 \$2011 \$1582 \$2010 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$928 \$2012 \$1582 \$2011 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$929 \$2013 \$1582 \$2012 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$930 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$931 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$932 \$2154 \$1581 \$1591 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$933 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$934 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$935 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$936 \$2156 \$1581 \$2155 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$937 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$938 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$939 \$2157 \$1581 \$1596 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$940 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$941 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$942 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$943 \$2159 \$1581 \$2158 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$944 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$945 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$946 \$2160 \$1581 \$1601 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$947 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$948 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$949 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$950 \$2161 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$951 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$952 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$953 \$2162 \$1582 \$1606 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$954 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$955 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$956 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$957 \$2163 \$1582 \$1611 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$958 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$959 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$960 \$2164 \$1582 \$1612 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$961 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$962 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$963 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$964 \$2165 \$1582 \$1617 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$965 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$966 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$967 \$2166 \$1582 \$1618 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$968 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$969 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$970 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$971 \$2167 \$1582 \$1623 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$972 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$973 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$974 \$2154 \$1581 \$2453 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$975 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$976 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$977 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$978 \$2156 \$1581 \$2454 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$979 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$980 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$981 \$2157 \$1581 \$2455 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$982 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$983 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$984 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$985 \$2159 \$1581 \$2456 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$986 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$987 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$988 \$2160 \$1581 \$2457 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$989 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$990 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$991 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$992 \$2161 \$1581 \$2458 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$993 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$994 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$995 \$2162 \$1582 \$2459 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$996 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$997 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$998 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$999 \$2163 \$1582 \$39 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1000 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1001 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1002 \$2164 \$1582 \$2460 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1003 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1004 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1005 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1006 \$2165 \$1582 \$40 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1007 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1008 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1009 \$2166 \$1582 \$2461 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1010 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1011 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1012 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1013 \$2167 \$1582 \$41 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1014 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1015 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1016 \$2718 \$1581 \$2717 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1017 \$2719 \$1581 \$2718 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1018 \$2720 \$1581 \$2719 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1019 \$2721 \$1581 \$2720 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1020 \$1988 \$1581 \$2721 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1021 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1022 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1023 \$2723 \$1581 \$2722 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1024 \$2724 \$1581 \$2723 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1025 \$2725 \$1581 \$2724 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1026 \$2726 \$1581 \$2725 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1027 \$1993 \$1581 \$2726 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1028 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1029 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1030 \$2728 \$1581 \$2727 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1031 \$2729 \$1581 \$2728 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1032 \$2730 \$1581 \$2729 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1033 \$2731 \$1581 \$2730 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1034 \$1998 \$1581 \$2731 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1035 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1036 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1037 \$2733 \$1582 \$2732 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1038 \$2734 \$1582 \$2733 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1039 \$2735 \$1582 \$2734 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1040 \$2736 \$1582 \$2735 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1041 \$2003 \$1582 \$2736 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1042 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1043 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1044 \$2738 \$1582 \$2737 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1045 \$2739 \$1582 \$2738 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1046 \$2740 \$1582 \$2739 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1047 \$2741 \$1582 \$2740 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1048 \$2008 \$1582 \$2741 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1049 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1050 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1051 \$2743 \$1582 \$2742 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1052 \$2744 \$1582 \$2743 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1053 \$2745 \$1582 \$2744 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1054 \$2746 \$1582 \$2745 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1055 \$2013 \$1582 \$2746 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1056 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1057 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1058 \$2961 \$1581 \$2717 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1059 \$2962 \$1581 \$2961 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1060 \$2963 \$1581 \$2962 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1061 \$2964 \$1581 \$2963 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1062 \$2965 \$1581 \$2964 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1063 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1064 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1065 \$2966 \$1581 \$2722 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1066 \$2967 \$1581 \$2966 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1067 \$2968 \$1581 \$2967 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1068 \$2969 \$1581 \$2968 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1069 \$2970 \$1581 \$2969 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1070 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1071 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1072 \$2971 \$1581 \$2727 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1073 \$2972 \$1581 \$2971 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1074 \$2973 \$1581 \$2972 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1075 \$2974 \$1581 \$2973 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1076 \$2975 \$1581 \$2974 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1077 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1078 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1079 \$2976 \$1582 \$2732 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1080 \$2977 \$1582 \$2976 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1081 \$2978 \$1582 \$2977 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1082 \$2979 \$1582 \$2978 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1083 \$2980 \$1582 \$2979 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1084 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1085 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1086 \$2981 \$1582 \$2737 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1087 \$2982 \$1582 \$2981 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1088 \$2983 \$1582 \$2982 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1089 \$2984 \$1582 \$2983 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1090 \$2985 \$1582 \$2984 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1091 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1092 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1093 \$2986 \$1582 \$2742 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1094 \$2987 \$1582 \$2986 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1095 \$2988 \$1582 \$2987 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1096 \$2989 \$1582 \$2988 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1097 \$2990 \$1582 \$2989 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1098 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1099 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1100 \$3273 \$1581 \$6536 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1101 \$3274 \$1581 \$3273 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1102 \$3275 \$1581 \$3274 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1103 \$3276 \$1581 \$3275 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1104 \$2965 \$1581 \$3276 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1105 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1106 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1107 \$3277 \$1581 \$6537 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1108 \$3278 \$1581 \$3277 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1109 \$3279 \$1581 \$3278 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1110 \$3280 \$1581 \$3279 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1111 \$2970 \$1581 \$3280 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1112 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1113 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1114 \$3282 \$1581 IBPOUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1115 \$3283 \$1581 \$3282 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1116 \$3284 \$1581 \$3283 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1117 \$3285 \$1581 \$3284 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1118 \$2975 \$1581 \$3285 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1119 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1120 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1121 \$3286 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1122 \$3287 \$1582 \$3286 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1123 \$3288 \$1582 \$3287 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1124 \$3289 \$1582 \$3288 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1125 \$2980 \$1582 \$3289 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1126 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1127 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1128 \$3290 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1129 \$3291 \$1582 \$3290 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1130 \$3292 \$1582 \$3291 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1131 \$3293 \$1582 \$3292 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1132 \$2985 \$1582 \$3293 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1133 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1134 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1135 \$3294 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1136 \$3295 \$1582 \$3294 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1137 \$3296 \$1582 \$3295 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1138 \$3297 \$1582 \$3296 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1139 \$2990 \$1582 \$3297 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1140 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1141 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1142 \$3541 \$1581 \$2453 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1143 \$3542 \$1581 \$3541 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1144 \$3543 \$1581 \$3542 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1145 \$3544 \$1581 \$3543 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1146 \$2454 \$1581 \$3544 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1147 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1148 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1149 \$3545 \$1581 \$2455 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1150 \$3546 \$1581 \$3545 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1151 \$3547 \$1581 \$3546 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1152 \$3548 \$1581 \$3547 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1153 \$2456 \$1581 \$3548 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1154 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1155 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1156 \$3549 \$1581 \$2457 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1157 \$3550 \$1581 \$3549 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1158 \$3551 \$1581 \$3550 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1159 \$3552 \$1581 \$3551 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1160 \$2458 \$1581 \$3552 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1161 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1162 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1163 \$3553 \$1582 \$2459 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1164 \$3554 \$1582 \$3553 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1165 \$3555 \$1582 \$3554 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1166 \$3556 \$1582 \$3555 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1167 VDD \$1582 \$3556 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1168 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1169 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1170 \$3557 \$1582 \$2460 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1171 \$3558 \$1582 \$3557 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1172 \$3559 \$1582 \$3558 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1173 \$3560 \$1582 \$3559 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1174 VDD \$1582 \$3560 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1175 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1176 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1177 \$3561 \$1582 \$2461 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1178 \$3562 \$1582 \$3561 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1179 \$3563 \$1582 \$3562 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1180 \$3564 \$1582 \$3563 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1181 VDD \$1582 \$3564 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1182 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1183 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1184 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1185 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1186 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1187 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1188 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1189 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1190 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1191 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1192 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1193 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1194 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1195 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1196 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1197 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1198 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1199 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1200 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1201 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1202 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1203 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1204 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1205 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1206 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1207 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1208 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1209 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1210 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1211 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1212 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1213 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1214 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1215 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1216 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1217 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1218 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1219 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1220 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1221 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1222 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1223 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1224 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1225 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1226 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1227 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1228 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1229 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1230 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1231 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1232 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1233 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1234 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1235 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1236 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1237 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1238 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1239 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1240 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1241 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1242 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1243 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1244 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1245 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1246 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1247 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1248 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1249 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1250 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1251 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1252 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1253 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1254 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1255 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1256 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1257 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1258 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1259 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1260 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1261 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1262 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1263 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1264 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1265 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1266 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1267 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1268 \$3880 \$1581 \$3879 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1269 \$3881 \$1581 \$3880 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1270 \$3882 \$1581 \$3881 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1271 \$3883 \$1581 \$3882 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1272 VDD \$1581 \$3883 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1273 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1274 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1275 \$3885 \$1581 \$3884 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1276 \$3886 \$1581 \$3885 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1277 \$3887 \$1581 \$3886 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1278 \$3888 \$1581 \$3887 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1279 VDD \$1581 \$3888 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1280 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1281 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1282 \$3890 \$1581 \$3889 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1283 \$3891 \$1581 \$3890 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1284 \$3892 \$1581 \$3891 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1285 \$3893 \$1581 \$3892 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1286 VDD \$1581 \$3893 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1287 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1288 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1289 \$3895 \$1582 \$3894 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1290 \$3896 \$1582 \$3895 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1291 \$3897 \$1582 \$3896 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1292 \$3898 \$1582 \$3897 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1293 \$3899 \$1582 \$3898 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1294 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1295 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1296 \$3901 \$1582 \$3900 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1297 \$3902 \$1582 \$3901 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1298 \$3903 \$1582 \$3902 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1299 \$3904 \$1582 \$3903 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1300 \$3905 \$1582 \$3904 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1301 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1302 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1303 \$3907 \$1582 \$3906 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1304 \$3908 \$1582 \$3907 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1305 \$3909 \$1582 \$3908 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1306 \$3910 \$1582 \$3909 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1307 \$3911 \$1582 \$3910 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1308 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1309 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1310 \$4054 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1311 \$4055 \$1581 \$4054 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1312 \$4056 \$1581 \$4055 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1313 \$4057 \$1581 \$4056 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1314 \$4058 \$1581 \$4057 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1315 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1316 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1317 \$4059 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1318 \$4060 \$1581 \$4059 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1319 \$4061 \$1581 \$4060 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1320 \$4062 \$1581 \$4061 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1321 \$4063 \$1581 \$4062 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1322 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1323 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1324 \$4064 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1325 \$4065 \$1581 \$4064 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1326 \$4066 \$1581 \$4065 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1327 \$4067 \$1581 \$4066 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1328 \$4068 \$1581 \$4067 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1329 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1330 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1331 \$4069 \$1582 \$187 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1332 \$4070 \$1582 \$4069 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1333 \$4071 \$1582 \$4070 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1334 \$4072 \$1582 \$4071 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1335 \$4073 \$1582 \$4072 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1336 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1337 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1338 \$4074 \$1582 \$189 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1339 \$4075 \$1582 \$4074 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1340 \$4076 \$1582 \$4075 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1341 \$4077 \$1582 \$4076 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1342 \$4078 \$1582 \$4077 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1343 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1344 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1345 \$4079 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1346 \$4080 \$1582 \$4079 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1347 \$4081 \$1582 \$4080 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1348 \$4082 \$1582 \$4081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1349 \$4083 \$1582 \$4082 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1350 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1351 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1352 \$4220 \$1581 \$4219 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1353 \$4221 \$1581 \$4220 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1354 \$4222 \$1581 \$4221 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1355 \$4223 \$1581 \$4222 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1356 \$4058 \$1581 \$4223 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1357 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1358 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1359 \$4225 \$1581 \$4224 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1360 \$4226 \$1581 \$4225 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1361 \$4227 \$1581 \$4226 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1362 \$4228 \$1581 \$4227 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1363 \$4063 \$1581 \$4228 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1364 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1365 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1366 \$4230 \$1581 \$4229 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1367 \$4231 \$1581 \$4230 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1368 \$4232 \$1581 \$4231 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1369 \$4233 \$1581 \$4232 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1370 \$4068 \$1581 \$4233 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1371 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1372 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1373 \$4235 \$1582 \$4234 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1374 \$4236 \$1582 \$4235 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1375 \$4237 \$1582 \$4236 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1376 \$4238 \$1582 \$4237 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1377 \$4073 \$1582 \$4238 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1378 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1379 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1380 \$4240 \$1582 \$4239 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1381 \$4241 \$1582 \$4240 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1382 \$4242 \$1582 \$4241 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1383 \$4243 \$1582 \$4242 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1384 \$4078 \$1582 \$4243 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1385 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1386 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1387 \$4245 \$1582 \$4244 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1388 \$4246 \$1582 \$4245 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1389 \$4247 \$1582 \$4246 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1390 \$4248 \$1582 \$4247 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1391 \$4083 \$1582 \$4248 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1392 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1393 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1394 \$4375 \$1581 \$4219 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1395 \$4376 \$1581 \$4375 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1396 \$4377 \$1581 \$4376 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1397 \$4378 \$1581 \$4377 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1398 \$4379 \$1581 \$4378 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1399 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1400 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1401 \$4380 \$1581 \$4224 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1402 \$4381 \$1581 \$4380 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1403 \$4382 \$1581 \$4381 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1404 \$4383 \$1581 \$4382 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1405 \$4384 \$1581 \$4383 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1406 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1407 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1408 \$4385 \$1581 \$4229 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1409 \$4386 \$1581 \$4385 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1410 \$4387 \$1581 \$4386 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1411 \$4388 \$1581 \$4387 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1412 \$4389 \$1581 \$4388 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1413 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1414 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1415 \$4390 \$1582 \$4234 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1416 \$4391 \$1582 \$4390 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1417 \$4392 \$1582 \$4391 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1418 \$4393 \$1582 \$4392 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1419 \$4394 \$1582 \$4393 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1420 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1421 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1422 \$4395 \$1582 \$4239 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1423 \$4396 \$1582 \$4395 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1424 \$4397 \$1582 \$4396 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1425 \$4398 \$1582 \$4397 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1426 \$4399 \$1582 \$4398 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1427 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1428 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1429 \$4400 \$1582 \$4244 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1430 \$4401 \$1582 \$4400 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1431 \$4402 \$1582 \$4401 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1432 \$4403 \$1582 \$4402 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1433 \$4404 \$1582 \$4403 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1434 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1435 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1436 \$4539 \$1581 \$3879 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1437 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1438 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1439 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1440 \$4540 \$1581 \$4557 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1441 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1442 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1443 \$4541 \$1581 \$3884 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1444 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1445 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1446 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1447 \$4542 \$1581 \$4558 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1448 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1449 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1450 \$4543 \$1581 \$3889 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1451 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1452 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1453 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1454 \$4544 \$1581 \$4559 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1455 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1456 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1457 \$4545 \$1582 \$3894 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1458 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1459 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1460 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1461 \$4546 \$1582 \$3899 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1462 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1463 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1464 \$4547 \$1582 \$3900 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1465 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1466 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1467 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1468 \$4548 \$1582 \$3905 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1469 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1470 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1471 \$4549 \$1582 \$3906 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1472 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1473 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1474 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1475 \$4550 \$1582 \$3911 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1476 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1477 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1478 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1479 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1480 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1481 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1482 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1483 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1484 \$4539 \$1581 \$4701 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1485 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1486 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1487 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1488 \$4540 \$1581 \$4702 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1489 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1490 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1491 \$4541 \$1581 \$4703 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1492 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1493 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1494 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1495 \$4542 \$1581 \$4704 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1496 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1497 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1498 \$4543 \$1581 \$4705 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1499 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1500 \$1581 \$1581 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1501 VDD \$1581 \$1581 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1502 \$4544 \$1581 \$4706 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1503 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1504 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1505 \$4545 \$1582 \$4707 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1506 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1507 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1508 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1509 \$4546 \$1582 \$42 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1510 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1511 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1512 \$4547 \$1582 \$4708 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1513 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1514 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1515 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1516 \$4548 \$1582 \$43 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1517 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1518 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1519 \$4549 \$1582 \$4709 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1520 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1521 VDD \$1582 \$1582 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1522 \$1582 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1523 \$4550 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1524 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1525 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1526 \$4742 \$4700 \$1769 VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1527 VDD \$4700 \$4742 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1528 \$4743 \$4700 VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1529 \$1770 \$4700 \$4743 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1530 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1531 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1532 \$4876 \$1581 \$4875 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1533 \$4877 \$1581 \$4876 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1534 \$4878 \$1581 \$4877 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1535 \$4879 \$1581 \$4878 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1536 \$4379 \$1581 \$4879 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1537 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1538 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1539 \$4881 \$1581 \$4880 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1540 \$4882 \$1581 \$4881 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1541 \$4883 \$1581 \$4882 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1542 \$4884 \$1581 \$4883 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1543 \$4384 \$1581 \$4884 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1544 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1545 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1546 \$4886 \$1581 \$4885 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1547 \$4887 \$1581 \$4886 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1548 \$4888 \$1581 \$4887 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1549 \$4889 \$1581 \$4888 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1550 \$4389 \$1581 \$4889 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1551 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1552 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1553 \$4891 \$1582 \$4890 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1554 \$4892 \$1582 \$4891 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1555 \$4893 \$1582 \$4892 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1556 \$4894 \$1582 \$4893 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1557 \$4394 \$1582 \$4894 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1558 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1559 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1560 \$4896 \$1582 \$4895 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1561 \$4897 \$1582 \$4896 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1562 \$4898 \$1582 \$4897 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1563 \$4899 \$1582 \$4898 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1564 \$4399 \$1582 \$4899 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1565 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1566 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1567 \$4901 \$1582 \$4900 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1568 \$4902 \$1582 \$4901 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1569 \$4903 \$1582 \$4902 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1570 \$4904 \$1582 \$4903 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1571 \$4404 \$1582 \$4904 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1572 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1573 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1574 \$4925 \$4700 \$4700 VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1575 VDD \$4700 \$4925 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1576 \$4926 \$4700 VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1577 \$4700 \$4700 \$4926 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1578 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1579 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1580 \$5064 \$1581 \$4875 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1581 \$5065 \$1581 \$5064 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1582 \$5066 \$1581 \$5065 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1583 \$5067 \$1581 \$5066 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1584 \$5068 \$1581 \$5067 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1585 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1586 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1587 \$5069 \$1581 \$4880 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1588 \$5070 \$1581 \$5069 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1589 \$5071 \$1581 \$5070 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1590 \$5072 \$1581 \$5071 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1591 \$5073 \$1581 \$5072 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1592 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1593 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1594 \$5074 \$1581 \$4885 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1595 \$5075 \$1581 \$5074 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1596 \$5076 \$1581 \$5075 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1597 \$5077 \$1581 \$5076 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1598 \$5078 \$1581 \$5077 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1599 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1600 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1601 \$5079 \$1582 \$4890 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1602 \$5080 \$1582 \$5079 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1603 \$5081 \$1582 \$5080 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1604 \$5082 \$1582 \$5081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1605 \$5083 \$1582 \$5082 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1606 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1607 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1608 \$5084 \$1582 \$4895 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1609 \$5085 \$1582 \$5084 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1610 \$5086 \$1582 \$5085 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1611 \$5087 \$1582 \$5086 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1612 \$5088 \$1582 \$5087 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1613 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1614 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1615 \$5089 \$1582 \$4900 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1616 \$5090 \$1582 \$5089 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1617 \$5091 \$1582 \$5090 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1618 \$5092 \$1582 \$5091 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1619 \$5093 \$1582 \$5092 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1620 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1621 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1622 \$5129 \$4700 \$1770 VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1623 VDD \$4700 \$5129 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1624 \$5130 \$4700 VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1625 \$1769 \$4700 \$5130 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1626 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1627 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1628 \$5222 \$1581 \$6533 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1629 \$5223 \$1581 \$5222 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1630 \$5224 \$1581 \$5223 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1631 \$5225 \$1581 \$5224 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1632 \$5068 \$1581 \$5225 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1633 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1634 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1635 \$5226 \$1581 \$6534 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1636 \$5227 \$1581 \$5226 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1637 \$5228 \$1581 \$5227 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1638 \$5229 \$1581 \$5228 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1639 \$5073 \$1581 \$5229 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1640 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1641 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1642 \$5230 \$1581 \$6535 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1643 \$5231 \$1581 \$5230 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1644 \$5232 \$1581 \$5231 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1645 \$5233 \$1581 \$5232 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1646 \$5078 \$1581 \$5233 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1647 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1648 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1649 \$5234 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1650 \$5235 \$1582 \$5234 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1651 \$5236 \$1582 \$5235 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1652 \$5237 \$1582 \$5236 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1653 \$5083 \$1582 \$5237 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1654 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1655 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1656 \$5238 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1657 \$5239 \$1582 \$5238 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1658 \$5240 \$1582 \$5239 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1659 \$5241 \$1582 \$5240 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1660 \$5088 \$1582 \$5241 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1661 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1662 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1663 \$5242 \$1582 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1664 \$5243 \$1582 \$5242 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1665 \$5244 \$1582 \$5243 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1666 \$5245 \$1582 \$5244 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1667 \$5093 \$1582 \$5245 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1668 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1669 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1670 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1671 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1672 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1673 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1674 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1675 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1676 \$5360 \$1581 \$4701 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1677 \$5361 \$1581 \$5360 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1678 \$5362 \$1581 \$5361 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1679 \$5363 \$1581 \$5362 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1680 \$4702 \$1581 \$5363 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1681 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1682 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1683 \$5364 \$1581 \$4703 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1684 \$5365 \$1581 \$5364 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1685 \$5366 \$1581 \$5365 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1686 \$5367 \$1581 \$5366 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1687 \$4704 \$1581 \$5367 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1688 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1689 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1690 \$5368 \$1581 \$4705 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1691 \$5369 \$1581 \$5368 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1692 \$5370 \$1581 \$5369 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1693 \$5371 \$1581 \$5370 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1694 \$4706 \$1581 \$5371 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1695 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1696 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1697 \$5372 \$1582 \$4707 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1698 \$5373 \$1582 \$5372 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1699 \$5374 \$1582 \$5373 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1700 \$5375 \$1582 \$5374 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1701 VDD \$1582 \$5375 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1702 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1703 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1704 \$5376 \$1582 \$4708 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1705 \$5377 \$1582 \$5376 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1706 \$5378 \$1582 \$5377 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1707 \$5379 \$1582 \$5378 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1708 VDD \$1582 \$5379 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1709 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1710 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1711 \$5380 \$1582 \$4709 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1712 \$5381 \$1582 \$5380 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1713 \$5382 \$1582 \$5381 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1714 \$5383 \$1582 \$5382 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1715 VDD \$1582 \$5383 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1716 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1717 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1718 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1719 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1720 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1721 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1722 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1723 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1724 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1725 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1726 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1727 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1728 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1729 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1730 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1731 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1732 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1733 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1734 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1735 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1736 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1737 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1738 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1739 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1740 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1741 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1742 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1743 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1744 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1745 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1746 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1747 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1748 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1749 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1750 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1751 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1752 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1753 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1754 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1755 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1756 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1757 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1758 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1759 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1760 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1761 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1762 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1763 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1764 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1765 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1766 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1767 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1768 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1769 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1770 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1771 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1772 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1773 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1774 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1775 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1776 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1777 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1778 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1779 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1780 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1781 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1782 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1783 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1784 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1785 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1786 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1787 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1788 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1789 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1790 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1791 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1792 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1793 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1794 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1795 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1796 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1797 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1798 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1799 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1800 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1801 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1802 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1803 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1804 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1805 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1806 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1807 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1808 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1809 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1810 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1811 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1812 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1813 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1814 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1815 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1816 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1817 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1818 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1819 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1820 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1821 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1822 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1823 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1824 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1825 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1826 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1827 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1828 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1829 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1830 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1831 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1832 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1833 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1834 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1835 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1836 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1837 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1838 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1839 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1840 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1841 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1842 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1843 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1844 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1845 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1846 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1847 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1848 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1849 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1850 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1851 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1852 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1853 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1854 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1855 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1856 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1857 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1858 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1859 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1860 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1861 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1862 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1863 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1864 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1865 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1866 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1867 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1868 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1869 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1870 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1871 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1872 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1873 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1874 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1875 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1876 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1877 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1878 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1879 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1880 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1881 \$6434 \$5689 \$5689 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1882 VDD \$5689 \$6434 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1883 \$6435 \$5689 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1884 \$5588 \$5689 \$6435 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1885 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1886 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1887 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1888 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1889 \$6436 \$6468 \$34238 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1890 \$5692 \$6468 \$6436 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1891 \$6437 \$6468 \$5799 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1892 \$6438 \$6468 \$6437 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1893 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1894 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1895 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1896 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1897 \$6439 \$5789 \$5790 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1898 \$4557 \$5789 \$6439 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1899 \$6440 \$6533 \$4557 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1900 \$6468 \$6533 \$6440 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1901 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1902 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1903 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1904 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1905 \$6441 \$5697 \$5697 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1906 VDD \$5697 \$6441 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1907 \$6442 \$5697 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1908 \$5589 \$5697 \$6442 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1909 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1910 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1911 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1912 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1913 \$6443 \$6469 \$6438 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1914 \$5700 \$6469 \$6443 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1915 \$6444 \$6469 \$5800 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1916 \$6445 \$6469 \$6444 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1917 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1918 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1919 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1920 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1921 \$6446 \$5791 \$5792 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1922 \$4558 \$5791 \$6446 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1923 \$6447 \$6534 \$4558 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1924 \$6469 \$6534 \$6447 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1925 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1926 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1927 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1928 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1929 \$6448 \$5705 \$5705 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1930 VDD \$5705 \$6448 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1931 \$6449 \$5705 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1932 \$5590 \$5705 \$6449 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1933 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1934 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1935 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1936 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1937 \$6450 \$6470 \$6445 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1938 \$5708 \$6470 \$6450 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1939 \$6451 \$6470 \$5801 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1940 \$6452 \$6470 \$6451 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1941 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1942 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1943 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1944 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1945 \$6453 \$5793 \$5794 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1946 \$4559 \$5793 \$6453 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1947 \$6454 \$6535 \$4559 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1948 \$6470 \$6535 \$6454 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1949 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1950 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1951 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1952 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1953 \$6455 \$5713 \$5713 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1954 VDD \$5713 \$6455 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1955 \$6456 \$5713 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1956 \$5591 \$5713 \$6456 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1957 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1958 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1959 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1960 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1961 \$6457 \$6471 \$6452 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1962 \$5716 \$6471 \$6457 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1963 \$6458 \$6471 \$5802 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1964 \$6459 \$6471 \$6458 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1965 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1966 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1967 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1968 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1969 \$6460 \$5795 \$5796 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1970 \$2155 \$5795 \$6460 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1971 \$6461 \$6536 \$2155 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1972 \$6471 \$6536 \$6461 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1973 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1974 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1975 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1976 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1977 \$6462 \$5721 \$5721 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1978 VDD \$5721 \$6462 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1979 \$6463 \$5721 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1980 \$5592 \$5721 \$6463 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1981 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1982 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1983 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1984 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1985 \$6464 \$6472 \$6459 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1986 \$5724 \$6472 \$6464 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1987 \$6465 \$6472 \$5803 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1988 OUT \$6472 \$6465 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1989 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1990 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1991 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1992 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1993 \$6466 \$5797 \$5798 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1994 \$2158 \$5797 \$6466 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1995 \$6467 \$6537 \$2158 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1996 \$6472 \$6537 \$6467 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1997 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1998 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1999 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2000 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2001 \$6608 \$5689 \$5588 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2002 VDD \$5689 \$6608 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2003 \$6609 \$5689 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2004 \$5689 \$5689 \$6609 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2005 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2006 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2007 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2008 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2009 \$6610 \$6468 \$6533 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2010 VSS \$6468 \$6610 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2011 \$6611 \$6468 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2012 \$6533 \$6468 \$6611 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2013 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2014 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2015 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2016 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2017 \$6612 \$6533 \$6468 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2018 \$4557 \$6533 \$6612 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2019 \$6613 \$5789 \$4557 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2020 \$5790 \$5789 \$6613 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2021 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2022 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2023 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2024 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2025 \$6614 \$5697 \$5589 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2026 VDD \$5697 \$6614 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2027 \$6615 \$5697 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2028 \$5697 \$5697 \$6615 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2029 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2030 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2031 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2032 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2033 \$6616 \$6469 \$6534 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2034 VSS \$6469 \$6616 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2035 \$6617 \$6469 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2036 \$6534 \$6469 \$6617 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2037 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2038 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2039 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2040 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2041 \$6618 \$6534 \$6469 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2042 \$4558 \$6534 \$6618 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2043 \$6619 \$5791 \$4558 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2044 \$5792 \$5791 \$6619 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2045 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2046 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2047 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2048 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2049 \$6620 \$5705 \$5590 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2050 VDD \$5705 \$6620 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2051 \$6621 \$5705 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2052 \$5705 \$5705 \$6621 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2053 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2054 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2055 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2056 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2057 \$6622 \$6470 \$6535 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2058 VSS \$6470 \$6622 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2059 \$6623 \$6470 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2060 \$6535 \$6470 \$6623 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2061 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2062 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2063 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2064 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2065 \$6624 \$6535 \$6470 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2066 \$4559 \$6535 \$6624 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2067 \$6625 \$5793 \$4559 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2068 \$5794 \$5793 \$6625 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2069 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2070 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2071 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2072 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2073 \$6626 \$5713 \$5591 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2074 VDD \$5713 \$6626 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2075 \$6627 \$5713 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2076 \$5713 \$5713 \$6627 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2077 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2078 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2079 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2080 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2081 \$6628 \$6471 \$6536 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2082 VSS \$6471 \$6628 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2083 \$6629 \$6471 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2084 \$6536 \$6471 \$6629 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2085 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2086 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2087 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2088 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2089 \$6630 \$6536 \$6471 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2090 \$2155 \$6536 \$6630 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2091 \$6631 \$5795 \$2155 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2092 \$5796 \$5795 \$6631 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2093 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2094 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2095 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2096 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2097 \$6632 \$5721 \$5592 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2098 VDD \$5721 \$6632 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2099 \$6633 \$5721 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2100 \$5721 \$5721 \$6633 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2101 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2102 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2103 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2104 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2105 \$6634 \$6472 \$6537 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2106 VSS \$6472 \$6634 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2107 \$6635 \$6472 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2108 \$6537 \$6472 \$6635 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2109 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2110 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2111 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2112 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2113 \$6636 \$6537 \$6472 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2114 \$2158 \$6537 \$6636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2115 \$6637 \$5797 \$2158 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2116 \$5798 \$5797 \$6637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2117 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2118 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2119 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2120 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2121 \$6729 \$5689 \$5689 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2122 VDD \$5689 \$6729 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2123 \$6730 \$5689 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2124 \$5588 \$5689 \$6730 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2125 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2126 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2127 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2128 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2129 \$6731 \$6468 \$6533 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2130 VSS \$6468 \$6731 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2131 \$6732 \$6468 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2132 \$6533 \$6468 \$6732 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2133 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2134 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2135 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2136 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2137 \$6733 \$5789 \$5790 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2138 \$4557 \$5789 \$6733 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2139 \$6734 \$6533 \$4557 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2140 \$6468 \$6533 \$6734 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2141 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2142 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2143 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2144 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2145 \$6735 \$5697 \$5697 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2146 VDD \$5697 \$6735 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2147 \$6736 \$5697 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2148 \$5589 \$5697 \$6736 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2149 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2150 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2151 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2152 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2153 \$6737 \$6469 \$6534 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2154 VSS \$6469 \$6737 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2155 \$6738 \$6469 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2156 \$6534 \$6469 \$6738 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2157 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2158 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2159 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2160 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2161 \$6739 \$5791 \$5792 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2162 \$4558 \$5791 \$6739 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2163 \$6740 \$6534 \$4558 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2164 \$6469 \$6534 \$6740 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2165 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2166 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2167 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2168 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2169 \$6741 \$5705 \$5705 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2170 VDD \$5705 \$6741 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2171 \$6742 \$5705 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2172 \$5590 \$5705 \$6742 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2173 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2174 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2175 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2176 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2177 \$6743 \$6470 \$6535 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2178 VSS \$6470 \$6743 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2179 \$6744 \$6470 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2180 \$6535 \$6470 \$6744 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2181 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2182 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2183 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2184 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2185 \$6745 \$5793 \$5794 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2186 \$4559 \$5793 \$6745 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2187 \$6746 \$6535 \$4559 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2188 \$6470 \$6535 \$6746 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2189 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2190 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2191 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2192 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2193 \$6747 \$5713 \$5713 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2194 VDD \$5713 \$6747 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2195 \$6748 \$5713 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2196 \$5591 \$5713 \$6748 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2197 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2198 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2199 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2200 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2201 \$6749 \$6471 \$6536 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2202 VSS \$6471 \$6749 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2203 \$6750 \$6471 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2204 \$6536 \$6471 \$6750 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2205 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2206 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2207 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2208 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2209 \$6751 \$5795 \$5796 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2210 \$2155 \$5795 \$6751 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2211 \$6752 \$6536 \$2155 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2212 \$6471 \$6536 \$6752 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2213 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2214 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2215 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2216 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2217 \$6753 \$5721 \$5721 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2218 VDD \$5721 \$6753 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2219 \$6754 \$5721 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2220 \$5592 \$5721 \$6754 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2221 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2222 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2223 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2224 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2225 \$6755 \$6472 \$6537 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2226 VSS \$6472 \$6755 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2227 \$6756 \$6472 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2228 \$6537 \$6472 \$6756 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2229 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2230 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2231 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2232 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2233 \$6757 \$5797 \$5798 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2234 \$2158 \$5797 \$6757 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2235 \$6758 \$6537 \$2158 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2236 \$6472 \$6537 \$6758 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2237 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2238 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2239 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2240 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2241 \$6874 \$5689 \$5588 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2242 VDD \$5689 \$6874 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2243 \$6875 \$5689 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2244 \$5689 \$5689 \$6875 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2245 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2246 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2247 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2248 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2249 \$6876 \$6468 \$6438 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2250 \$5799 \$6468 \$6876 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2251 \$6877 \$6468 \$5692 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2252 \$34238 \$6468 \$6877 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2253 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2254 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2255 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2256 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2257 \$6878 \$6533 \$6468 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2258 \$4557 \$6533 \$6878 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2259 \$6879 \$5789 \$4557 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2260 \$5790 \$5789 \$6879 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2261 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2262 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2263 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2264 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2265 \$6880 \$5697 \$5589 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2266 VDD \$5697 \$6880 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2267 \$6881 \$5697 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2268 \$5697 \$5697 \$6881 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2269 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2270 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2271 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2272 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2273 \$6882 \$6469 \$6445 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2274 \$5800 \$6469 \$6882 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2275 \$6883 \$6469 \$5700 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2276 \$6438 \$6469 \$6883 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2277 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2278 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2279 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2280 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2281 \$6884 \$6534 \$6469 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2282 \$4558 \$6534 \$6884 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2283 \$6885 \$5791 \$4558 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2284 \$5792 \$5791 \$6885 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2285 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2286 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2287 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2288 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2289 \$6886 \$5705 \$5590 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2290 VDD \$5705 \$6886 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2291 \$6887 \$5705 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2292 \$5705 \$5705 \$6887 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2293 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2294 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2295 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2296 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2297 \$6888 \$6470 \$6452 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2298 \$5801 \$6470 \$6888 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2299 \$6889 \$6470 \$5708 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2300 \$6445 \$6470 \$6889 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2301 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2302 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2303 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2304 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2305 \$6890 \$6535 \$6470 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2306 \$4559 \$6535 \$6890 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2307 \$6891 \$5793 \$4559 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2308 \$5794 \$5793 \$6891 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2309 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2310 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2311 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2312 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2313 \$6892 \$5713 \$5591 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2314 VDD \$5713 \$6892 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2315 \$6893 \$5713 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2316 \$5713 \$5713 \$6893 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2317 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2318 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2319 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2320 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2321 \$6894 \$6471 \$6459 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2322 \$5802 \$6471 \$6894 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2323 \$6895 \$6471 \$5716 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2324 \$6452 \$6471 \$6895 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2325 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2326 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2327 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2328 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2329 \$6896 \$6536 \$6471 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2330 \$2155 \$6536 \$6896 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2331 \$6897 \$5795 \$2155 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2332 \$5796 \$5795 \$6897 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2333 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2334 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2335 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2336 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2337 \$6898 \$5721 \$5592 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2338 VDD \$5721 \$6898 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2339 \$6899 \$5721 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2340 \$5721 \$5721 \$6899 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2341 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2342 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2343 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2344 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2345 \$6900 \$6472 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2346 \$5803 \$6472 \$6900 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2347 \$6901 \$6472 \$5724 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2348 \$6459 \$6472 \$6901 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2349 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2350 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2351 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2352 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2353 \$6902 \$6537 \$6472 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2354 \$2158 \$6537 \$6902 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2355 \$6903 \$5797 \$2158 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2356 \$5798 \$5797 \$6903 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2357 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2358 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2359 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2360 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2361 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2362 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2363 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2364 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2365 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2366 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2367 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2368 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2369 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2370 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2371 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2372 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2373 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2374 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2375 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2376 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2377 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2378 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2379 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2380 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2381 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2382 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2383 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2384 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2385 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2386 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2387 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2388 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2389 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2390 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2391 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2392 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2393 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2394 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2395 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2396 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2397 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2398 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2399 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2400 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2401 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2402 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2403 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2404 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2405 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2406 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2407 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2408 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2409 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2410 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2411 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2412 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2413 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2414 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2415 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2416 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2417 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2418 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2419 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2420 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2421 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2422 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2423 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2424 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2425 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2426 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2427 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2428 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2429 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2430 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2431 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2432 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2433 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2434 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2435 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2436 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2437 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2438 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2439 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2440 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2441 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2442 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2443 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2444 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2445 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2446 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2447 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2448 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2449 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2450 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2451 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2452 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2453 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2454 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2455 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2456 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2457 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2458 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2459 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2460 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2461 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2462 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2463 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2464 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2465 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2466 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2467 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2468 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2469 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2470 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2471 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2472 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2473 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2474 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2475 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2476 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2477 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2478 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2479 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2480 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2481 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2482 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2483 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2484 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2485 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2486 VDD \$10111 \$7132 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2487 \$7132 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2488 VDD \$10111 \$7132 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2489 \$7132 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2490 VDD \$10111 \$7693 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2491 \$7693 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2492 VDD \$10111 \$7693 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2493 \$7693 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2494 VDD \$10111 \$10111 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2495 \$10111 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2496 VDD \$10111 \$10111 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2497 \$10111 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2498 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2499 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2500 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2501 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2502 VDD \$10111 \$10111 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2503 \$10111 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2504 VDD \$10111 \$10111 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2505 \$10111 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2506 VDD \$10111 \$7693 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2507 \$7693 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2508 VDD \$10111 \$7693 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2509 \$7693 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2510 VDD \$10111 \$7132 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2511 \$7132 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2512 VDD \$10111 \$7132 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2513 \$7132 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2514 VDD \$10111 \$10111 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2515 \$10111 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2516 VDD \$10111 \$10111 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2517 VDD \$10111 \$7693 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2518 \$7693 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2519 VDD \$10111 \$7693 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2520 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2521 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2522 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2523 \$7693 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2524 VDD \$10111 \$7693 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2525 \$7693 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2526 \$7132 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2527 VDD \$10111 \$7132 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2528 \$7132 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2529 VDD \$10111 \$7132 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2530 \$7132 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2531 VDD \$10111 \$7132 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2532 VDD \$10111 \$10111 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2533 \$10111 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2534 VDD \$10111 \$10111 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2535 VDD \$10111 \$10111 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2536 \$10111 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2537 VDD \$10111 \$10111 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2538 \$10111 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2539 VDD \$10111 \$7693 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2540 \$7693 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2541 VDD \$10111 \$7693 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2542 \$7693 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2543 VDD \$10111 \$7693 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2544 \$7693 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2545 VDD \$10111 \$7693 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2546 \$7693 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2547 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2548 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2549 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2550 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2551 VDD \$10111 \$7132 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2552 \$7132 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2553 VDD \$10111 \$7132 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2554 \$7132 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2555 VDD \$10111 \$10111 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2556 \$10111 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2557 VDD \$10111 \$10111 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2558 \$10111 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2559 VDD \$10111 \$7132 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2560 \$7132 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2561 VDD \$10111 \$7132 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2562 \$7132 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2563 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2564 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2565 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2566 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2567 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2568 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2569 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2570 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2571 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2572 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2573 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2574 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2575 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2576 \$14901 \$7118 \$13568 VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P
+ PS=3.7U PD=2.04U
M$2577 \$14902 \$7118 \$14901 VDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P
+ PS=2.04U PD=2.04U
M$2578 \$14903 \$7118 \$14902 VDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P
+ PS=2.04U PD=3.7U
M$2579 \$15967 \$7118 \$15966 VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P
+ PS=3.7U PD=2.04U
M$2580 \$15968 \$7118 \$15967 VDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P
+ PS=2.04U PD=2.04U
M$2581 \$14903 \$7118 \$15968 VDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P
+ PS=2.04U PD=3.7U
M$2582 \$13569 \$7118 \$13568 VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P
+ PS=3.7U PD=2.04U
M$2583 \$13570 \$7118 \$13569 VDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P
+ PS=2.04U PD=2.04U
M$2584 VDD \$7118 \$13570 VDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P PS=2.04U
+ PD=3.7U
M$2585 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P PS=3.7U PD=2.04U
M$2586 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P PS=2.04U
+ PD=2.04U
M$2587 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P PS=2.04U PD=3.7U
M$2588 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P PS=3.7U PD=2.04U
M$2589 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P PS=2.04U
+ PD=2.04U
M$2590 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P PS=2.04U PD=3.7U
M$2591 \$17027 \$7118 \$15966 VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P
+ PS=3.7U PD=2.04U
M$2592 \$17028 \$7118 \$17027 VDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P
+ PS=2.04U PD=2.04U
M$2593 \$17029 \$7118 \$17028 VDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P
+ PS=2.04U PD=3.7U
M$2594 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2595 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2596 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2597 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2598 \$7118 \$7118 \$17029 VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P
+ PS=3.7U PD=3.7U
M$2599 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2600 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2601 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2602 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2603 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2604 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2605 VDD VDD VDD VDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$2606 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2607 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2608 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2609 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2610 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2611 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2612 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2613 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2614 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2615 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2616 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2617 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2618 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2619 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2620 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2621 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2622 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2623 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2624 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2625 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2626 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2627 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2628 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2629 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2630 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2631 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2632 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2633 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2634 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2635 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2636 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2637 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2638 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2639 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2640 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2641 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2642 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2643 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2644 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2645 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2646 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2647 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2648 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2649 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2650 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2651 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2652 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2653 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2654 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2655 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2656 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2657 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2658 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2659 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2660 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2661 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2662 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2663 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2664 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2665 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2666 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2667 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2668 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2669 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2670 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2671 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2672 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2673 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2674 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2675 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2676 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2677 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2678 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2679 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2680 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2681 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2682 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2683 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2684 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2685 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2686 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2687 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2688 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2689 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2690 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2691 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2692 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2693 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2694 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2695 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2696 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2697 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2698 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2699 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2700 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2701 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2702 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2703 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2704 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2705 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2706 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2707 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2708 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2709 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2710 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2711 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2712 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2713 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2714 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2715 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2716 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2717 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2718 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2719 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2720 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2721 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2722 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2723 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2724 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2725 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2726 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2727 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2728 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2729 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2730 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2731 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2732 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2733 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2734 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2735 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2736 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2737 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2738 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2739 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2740 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2741 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2742 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2743 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2744 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2745 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2746 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2747 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2748 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2749 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2750 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2751 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2752 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2753 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2754 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2755 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2756 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2757 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2758 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2759 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2760 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2761 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2762 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2763 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2764 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2765 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2766 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2767 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2768 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2769 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2770 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2771 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2772 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2773 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2774 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2775 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2776 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2777 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2778 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2779 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2780 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2781 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2782 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2783 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2784 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2785 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2786 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2787 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2788 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2789 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2790 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2791 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2792 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2793 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2794 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2795 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2796 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2797 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2798 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2799 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2800 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2801 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2802 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2803 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2804 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2805 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2806 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2807 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2808 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2809 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2810 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2811 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2812 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2813 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2814 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2815 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2816 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2817 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2818 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2819 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2820 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2821 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2822 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2823 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2824 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2825 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2826 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2827 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2828 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2829 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2830 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2831 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2832 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2833 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2834 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2835 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2836 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2837 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2838 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2839 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2840 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2841 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2842 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2843 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2844 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2845 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2846 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2847 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2848 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2849 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2850 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2851 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2852 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2853 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2854 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2855 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2856 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2857 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2858 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2859 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2860 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2861 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2862 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2863 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2864 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2865 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2866 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2867 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2868 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2869 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2870 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2871 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2872 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2873 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2874 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2875 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2876 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2877 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2878 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2879 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2880 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2881 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2882 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2883 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2884 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2885 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2886 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2887 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2888 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2889 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2890 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2891 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2892 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2893 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2894 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2895 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2896 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2897 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2898 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2899 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2900 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2901 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2902 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2903 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2904 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2905 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2906 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2907 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2908 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2909 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2910 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2911 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2912 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2913 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2914 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2915 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2916 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2917 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2918 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2919 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2920 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2921 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2922 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2923 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2924 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2925 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2926 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2927 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2928 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2929 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2930 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2931 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2932 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2933 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2934 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2935 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2936 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2937 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2938 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2939 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2940 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2941 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2942 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2943 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2944 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2945 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2946 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2947 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2948 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2949 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2950 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2951 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2952 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2953 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2954 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2955 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2956 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2957 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2958 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2959 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2960 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2961 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2962 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2963 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2964 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2965 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2966 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2967 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2968 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2969 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2970 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2971 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2972 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2973 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2974 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2975 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2976 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2977 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2978 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2979 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2980 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$2981 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2982 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2983 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2984 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2985 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2986 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2987 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2988 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2989 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2990 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2991 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2992 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2993 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2994 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2995 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2996 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2997 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2998 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2999 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3000 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3001 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3002 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3003 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3004 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3005 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3006 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3007 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3008 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3009 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3010 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3011 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3012 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3013 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3014 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3015 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3016 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3017 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3018 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3019 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3020 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3021 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3022 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3023 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3024 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3025 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3026 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3027 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3028 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3029 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3030 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3031 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3032 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3033 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3034 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3035 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3036 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3037 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3038 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3039 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3040 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3041 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3042 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3043 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3044 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3045 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3046 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3047 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3048 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3049 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3050 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3051 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3052 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3053 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3054 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3055 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3056 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3057 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3058 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3059 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3060 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3061 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3062 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3063 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3064 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3065 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3066 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3067 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3068 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3069 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3070 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3071 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3072 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3073 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3074 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3075 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3076 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3077 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3078 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3079 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3080 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3081 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3082 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3083 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3084 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3085 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3086 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3087 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3088 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3089 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3090 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3091 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3092 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3093 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3094 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3095 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3096 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3097 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3098 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3099 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3100 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3101 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3102 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3103 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3104 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3105 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3106 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3107 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3108 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3109 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3110 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3111 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3112 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3113 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3114 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3115 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3116 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3117 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3118 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3119 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3120 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3121 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3122 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3123 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3124 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3125 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3126 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3127 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3128 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3129 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3130 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3131 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3132 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3133 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3134 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3135 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3136 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3137 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3138 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3139 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3140 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3141 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3142 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3143 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3144 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3145 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3146 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3147 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3148 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3149 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3150 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3151 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3152 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3153 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3154 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3155 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3156 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3157 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3158 \$32636 \$34238 \$7081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3159 \$7081 \$34238 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3160 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3161 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3162 \$32636 \$6 \$7113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3163 \$7113 \$6 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3164 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3165 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3166 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3167 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3168 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3169 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3170 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3171 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3172 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3173 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3174 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3175 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3176 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3177 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3178 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3179 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3180 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3181 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3182 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3183 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3184 \$32638 \$7118 OUT VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3185 OUT \$7118 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3186 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3187 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3188 \$32637 \$7118 \$17566 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3189 \$17566 \$7118 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3190 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3191 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3192 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3193 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3194 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3195 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3196 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3197 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3198 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3199 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3200 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3201 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3202 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3203 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3204 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3205 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3206 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3207 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3208 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3209 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3210 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3211 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3212 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3213 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3214 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3215 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3216 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3217 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3218 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3219 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3220 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3221 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3222 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3223 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3224 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3225 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3226 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3227 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3228 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3229 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3230 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3231 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3232 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3233 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3234 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3235 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3236 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3237 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3238 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3239 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3240 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3241 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3242 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3243 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3244 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3245 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3246 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3247 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3248 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3249 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3250 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3251 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3252 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3253 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3254 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3255 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3256 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3257 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3258 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3259 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3260 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3261 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3262 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3263 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3264 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3265 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3266 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3267 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3268 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3269 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3270 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3271 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3272 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3273 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3274 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3275 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3276 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3277 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3278 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3279 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3280 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3281 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3282 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3283 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3284 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3285 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3286 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3287 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3288 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3289 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3290 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3291 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3292 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3293 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3294 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3295 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3296 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3297 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3298 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3299 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3300 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3301 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3302 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3303 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3304 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3305 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3306 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3307 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3308 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3309 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3310 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3311 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3312 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3313 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3314 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3315 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3316 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3317 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3318 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3319 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3320 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3321 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3322 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3323 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3324 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3325 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3326 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3327 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3328 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3329 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3330 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3331 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3332 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3333 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3334 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3335 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3336 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3337 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3338 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3339 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3340 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3341 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3342 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3343 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3344 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3345 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3346 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3347 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3348 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3349 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3350 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3351 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3352 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3353 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3354 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3355 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3356 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3357 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3358 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3359 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3360 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3361 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3362 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3363 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3364 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3365 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3366 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3367 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3368 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3369 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3370 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3371 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3372 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3373 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3374 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3375 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3376 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3377 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3378 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3379 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3380 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3381 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3382 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3383 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3384 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3385 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3386 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3387 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3388 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3389 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3390 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3391 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3392 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3393 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3394 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3395 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3396 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3397 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3398 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3399 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3400 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3401 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3402 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3403 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3404 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3405 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3406 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3407 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3408 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3409 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3410 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3411 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3412 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3413 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3414 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3415 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3416 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3417 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3418 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3419 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3420 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3421 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3422 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3423 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3424 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3425 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3426 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3427 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3428 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3429 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3430 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3431 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3432 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3433 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3434 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3435 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3436 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3437 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3438 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3439 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3440 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3441 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3442 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3443 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3444 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3445 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3446 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3447 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3448 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3449 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3450 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3451 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3452 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3453 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3454 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3455 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3456 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3457 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3458 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3459 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3460 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3461 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3462 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3463 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3464 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3465 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3466 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3467 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3468 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3469 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3470 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3471 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3472 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3473 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3474 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3475 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3476 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3477 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3478 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3479 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3480 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3481 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3482 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3483 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3484 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3485 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3486 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3487 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3488 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3489 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3490 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3491 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3492 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3493 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3494 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3495 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3496 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3497 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3498 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3499 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3500 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3501 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3502 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3503 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3504 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3505 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3506 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3507 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3508 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3509 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3510 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3511 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3512 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3513 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3514 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3515 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3516 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3517 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3518 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3519 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3520 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3521 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3522 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3523 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3524 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3525 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3526 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3527 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3528 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3529 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3530 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3531 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3532 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3533 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3534 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3535 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3536 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3537 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3538 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3539 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3540 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3541 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3542 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3543 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3544 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3545 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3546 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3547 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3548 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3549 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3550 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3551 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3552 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3553 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3554 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3555 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3556 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3557 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3558 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3559 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3560 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3561 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3562 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3563 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3564 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3565 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3566 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3567 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3568 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3569 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3570 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3571 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3572 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3573 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3574 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3575 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3576 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3577 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3578 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3579 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3580 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3581 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3582 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3583 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3584 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3585 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3586 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3587 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3588 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3589 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3590 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3591 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3592 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3593 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3594 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3595 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3596 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3597 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3598 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3599 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3600 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3601 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3602 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3603 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3604 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3605 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3606 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3607 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3608 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3609 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3610 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3611 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3612 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3613 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3614 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3615 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3616 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3617 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3618 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3619 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3620 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3621 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3622 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3623 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3624 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3625 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3626 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3627 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3628 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3629 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3630 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3631 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3632 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3633 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3634 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3635 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3636 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3637 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3638 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3639 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3640 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3641 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3642 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3643 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3644 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3645 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3646 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3647 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3648 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3649 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3650 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3651 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3652 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3653 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3654 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3655 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3656 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3657 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3658 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3659 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3660 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3661 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3662 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3663 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3664 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3665 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3666 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3667 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3668 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3669 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3670 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3671 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3672 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3673 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3674 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3675 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3676 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3677 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3678 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3679 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3680 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3681 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3682 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3683 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3684 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3685 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3686 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3687 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3688 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3689 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3690 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3691 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3692 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3693 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3694 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3695 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3696 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3697 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3698 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3699 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3700 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3701 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3702 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3703 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3704 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3705 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3706 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3707 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3708 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3709 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3710 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3711 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3712 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3713 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3714 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3715 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3716 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3717 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3718 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3719 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3720 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3721 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3722 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3723 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3724 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3725 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3726 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3727 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3728 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3729 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3730 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3731 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3732 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3733 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3734 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3735 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3736 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3737 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3738 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3739 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3740 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3741 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3742 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3743 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3744 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3745 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3746 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3747 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3748 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3749 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3750 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3751 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3752 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3753 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3754 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3755 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3756 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3757 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3758 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3759 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3760 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3761 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3762 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3763 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3764 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3765 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3766 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3767 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3768 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3769 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3770 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3771 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3772 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3773 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3774 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3775 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3776 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3777 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3778 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3779 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3780 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3781 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3782 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3783 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3784 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3785 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3786 VDD \$10111 \$32636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3787 \$32636 \$10111 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3788 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3789 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3790 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3791 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3792 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3793 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3794 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3795 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3796 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3797 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3798 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3799 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3800 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3801 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3802 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3803 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3804 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3805 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3806 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3807 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3808 VDD \$17566 \$32638 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3809 \$32638 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3810 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3811 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3812 VDD \$17566 \$32637 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3813 \$32637 \$17566 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3814 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3815 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3816 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3817 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3818 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3819 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3820 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3821 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3822 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3823 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3824 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3825 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3826 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3827 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3828 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3829 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3830 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3831 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3832 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3833 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3834 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3835 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3836 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3837 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3838 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3839 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3840 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3841 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3842 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3843 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3844 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3845 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3846 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3847 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3848 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3849 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3850 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3851 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3852 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3853 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3854 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3855 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3856 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3857 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3858 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3859 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3860 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3861 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3862 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3863 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3864 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$3865 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3866 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3867 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3868 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3869 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3870 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3871 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3872 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3873 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3874 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3875 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3876 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3877 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3878 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3879 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3880 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3881 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3882 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3883 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3884 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3885 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3886 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3887 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3888 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3889 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3890 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3891 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3892 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3893 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3894 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3895 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3896 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3897 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3898 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3899 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3900 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3901 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3902 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3903 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3904 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3905 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3906 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3907 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3908 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3909 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3910 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3911 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3912 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3913 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3914 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3915 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3916 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3917 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3918 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3919 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3920 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3921 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3922 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3923 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3924 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3925 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3926 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3927 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3928 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3929 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3930 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3931 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3932 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3933 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3934 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3935 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3936 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3937 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3938 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3939 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3940 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3941 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3942 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3943 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3944 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3945 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3946 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3947 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3948 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3949 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3950 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3951 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3952 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3953 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3954 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3955 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3956 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3957 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3958 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3959 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3960 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3961 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3962 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3963 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3964 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3965 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3966 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3967 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3968 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3969 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3970 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3971 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3972 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3973 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3974 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3975 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3976 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3977 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3978 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3979 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3980 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3981 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3982 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3983 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3984 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3985 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3986 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3987 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3988 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3989 \$894 \$924 \$925 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$3990 \$874 \$924 \$894 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$3991 \$895 \$266 \$874 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$3992 \$180 \$266 \$895 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$3993 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3994 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3995 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3996 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3997 \$896 \$925 \$148 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$3998 \$266 \$925 \$896 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$3999 \$897 \$925 \$266 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4000 \$125 \$925 \$897 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4001 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4002 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4003 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4004 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4005 \$898 \$265 \$34 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4006 VSS \$265 \$898 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4007 \$899 \$265 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4008 \$265 \$265 \$899 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4009 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4010 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4011 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4012 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4013 \$900 \$926 \$927 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4014 \$875 \$926 \$900 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4015 \$901 \$268 \$875 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4016 \$182 \$268 \$901 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4017 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4018 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4019 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4020 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4021 \$902 \$927 \$155 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4022 \$268 \$927 \$902 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4023 \$903 \$927 \$268 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4024 \$126 \$927 \$903 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4025 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4026 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4027 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4028 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4029 \$904 \$267 \$35 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4030 VSS \$267 \$904 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4031 \$905 \$267 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4032 \$267 \$267 \$905 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4033 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4034 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4035 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4036 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4037 \$906 \$928 \$929 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4038 \$876 \$928 \$906 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4039 \$907 \$270 \$876 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4040 \$184 \$270 \$907 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4041 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4042 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4043 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4044 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4045 \$908 \$929 \$162 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4046 \$270 \$929 \$908 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4047 \$909 \$929 \$270 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4048 \$127 \$929 \$909 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4049 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4050 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4051 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4052 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4053 \$910 \$269 \$36 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4054 VSS \$269 \$910 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4055 \$911 \$269 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4056 \$269 \$269 \$911 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4057 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4058 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4059 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4060 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4061 \$912 \$930 \$931 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4062 \$877 \$930 \$912 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4063 \$913 \$272 \$877 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4064 \$186 \$272 \$913 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4065 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4066 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4067 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4068 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4069 \$914 \$931 \$169 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4070 \$272 \$931 \$914 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4071 \$915 \$931 \$272 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4072 \$128 \$931 \$915 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4073 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4074 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4075 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4076 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4077 \$916 \$271 \$37 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4078 VSS \$271 \$916 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4079 \$917 \$271 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4080 \$271 \$271 \$917 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4081 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4082 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4083 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4084 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4085 \$918 \$932 \$933 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4086 \$878 \$932 \$918 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4087 \$919 \$274 \$878 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4088 \$188 \$274 \$919 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4089 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4090 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4091 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4092 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4093 \$920 \$933 \$176 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4094 \$274 \$933 \$920 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4095 \$921 \$933 \$274 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4096 \$129 \$933 \$921 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4097 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4098 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4099 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4100 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4101 \$922 \$273 \$38 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4102 VSS \$273 \$922 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4103 \$923 \$273 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4104 \$273 \$273 \$923 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4105 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4106 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4107 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4108 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4109 \$1049 \$266 \$180 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4110 \$874 \$266 \$1049 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4111 \$1050 \$924 \$874 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4112 \$925 \$924 \$1050 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4113 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4114 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4115 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4116 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4117 \$1051 \$925 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4118 \$924 \$925 \$1051 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4119 \$1052 \$925 \$924 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4120 VDD \$925 \$1052 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4121 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4122 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4123 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4124 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4125 \$1053 \$265 \$265 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4126 VSS \$265 \$1053 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4127 \$1054 \$265 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4128 \$34 \$265 \$1054 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4129 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4130 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4131 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4132 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4133 \$1055 \$268 \$182 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4134 \$875 \$268 \$1055 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4135 \$1056 \$926 \$875 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4136 \$927 \$926 \$1056 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4137 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4138 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4139 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4140 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4141 \$1057 \$927 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4142 \$926 \$927 \$1057 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4143 \$1058 \$927 \$926 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4144 VDD \$927 \$1058 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4145 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4146 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4147 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4148 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4149 \$1059 \$267 \$267 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4150 VSS \$267 \$1059 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4151 \$1060 \$267 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4152 \$35 \$267 \$1060 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4153 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4154 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4155 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4156 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4157 \$1061 \$270 \$184 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4158 \$876 \$270 \$1061 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4159 \$1062 \$928 \$876 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4160 \$929 \$928 \$1062 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4161 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4162 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4163 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4164 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4165 \$1063 \$929 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4166 \$928 \$929 \$1063 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4167 \$1064 \$929 \$928 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4168 VDD \$929 \$1064 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4169 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4170 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4171 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4172 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4173 \$1065 \$269 \$269 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4174 VSS \$269 \$1065 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4175 \$1066 \$269 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4176 \$36 \$269 \$1066 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4177 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4178 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4179 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4180 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4181 \$1067 \$272 \$186 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4182 \$877 \$272 \$1067 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4183 \$1068 \$930 \$877 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4184 \$931 \$930 \$1068 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4185 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4186 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4187 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4188 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4189 \$1069 \$931 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4190 \$930 \$931 \$1069 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4191 \$1070 \$931 \$930 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4192 VDD \$931 \$1070 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4193 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4194 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4195 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4196 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4197 \$1071 \$271 \$271 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4198 VSS \$271 \$1071 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4199 \$1072 \$271 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4200 \$37 \$271 \$1072 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4201 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4202 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4203 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4204 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4205 \$1073 \$274 \$188 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4206 \$878 \$274 \$1073 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4207 \$1074 \$932 \$878 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4208 \$933 \$932 \$1074 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4209 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4210 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4211 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4212 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4213 \$1075 \$933 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4214 \$932 \$933 \$1075 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4215 \$1076 \$933 \$932 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4216 VDD \$933 \$1076 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4217 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4218 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4219 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4220 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4221 \$1077 \$273 \$273 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4222 VSS \$273 \$1077 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4223 \$1078 \$273 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4224 \$38 \$273 \$1078 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4225 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4226 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4227 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4228 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4229 \$1184 \$924 \$925 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4230 \$874 \$924 \$1184 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4231 \$1185 \$266 \$874 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4232 \$180 \$266 \$1185 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4233 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4234 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4235 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4236 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4237 \$1186 \$925 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4238 \$924 \$925 \$1186 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4239 \$1187 \$925 \$924 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4240 VDD \$925 \$1187 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4241 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4242 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4243 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4244 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4245 \$1188 \$265 \$34 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4246 VSS \$265 \$1188 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4247 \$1189 \$265 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4248 \$265 \$265 \$1189 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4249 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4250 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4251 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4252 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4253 \$1190 \$926 \$927 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4254 \$875 \$926 \$1190 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4255 \$1191 \$268 \$875 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4256 \$182 \$268 \$1191 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4257 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4258 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4259 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4260 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4261 \$1192 \$927 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4262 \$926 \$927 \$1192 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4263 \$1193 \$927 \$926 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4264 VDD \$927 \$1193 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4265 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4266 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4267 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4268 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4269 \$1194 \$267 \$35 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4270 VSS \$267 \$1194 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4271 \$1195 \$267 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4272 \$267 \$267 \$1195 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4273 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4274 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4275 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4276 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4277 \$1196 \$928 \$929 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4278 \$876 \$928 \$1196 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4279 \$1197 \$270 \$876 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4280 \$184 \$270 \$1197 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4281 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4282 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4283 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4284 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4285 \$1198 \$929 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4286 \$928 \$929 \$1198 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4287 \$1199 \$929 \$928 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4288 VDD \$929 \$1199 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4289 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4290 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4291 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4292 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4293 \$1200 \$269 \$36 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4294 VSS \$269 \$1200 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4295 \$1201 \$269 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4296 \$269 \$269 \$1201 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4297 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4298 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4299 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4300 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4301 \$1202 \$930 \$931 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4302 \$877 \$930 \$1202 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4303 \$1203 \$272 \$877 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4304 \$186 \$272 \$1203 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4305 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4306 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4307 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4308 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4309 \$1204 \$931 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4310 \$930 \$931 \$1204 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4311 \$1205 \$931 \$930 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4312 VDD \$931 \$1205 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4313 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4314 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4315 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4316 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4317 \$1206 \$271 \$37 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4318 VSS \$271 \$1206 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4319 \$1207 \$271 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4320 \$271 \$271 \$1207 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4321 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4322 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4323 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4324 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4325 \$1208 \$932 \$933 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4326 \$878 \$932 \$1208 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4327 \$1209 \$274 \$878 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4328 \$188 \$274 \$1209 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4329 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4330 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4331 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4332 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4333 \$1210 \$933 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4334 \$932 \$933 \$1210 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4335 \$1211 \$933 \$932 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4336 VDD \$933 \$1211 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4337 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4338 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4339 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4340 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4341 \$1212 \$273 \$38 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4342 VSS \$273 \$1212 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4343 \$1213 \$273 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4344 \$273 \$273 \$1213 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4345 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4346 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4347 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4348 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4349 \$1329 \$266 \$180 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4350 \$874 \$266 \$1329 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4351 \$1330 \$924 \$874 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4352 \$925 \$924 \$1330 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4353 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4354 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4355 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4356 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4357 \$1331 \$925 \$125 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4358 \$266 \$925 \$1331 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4359 \$1332 \$925 \$266 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4360 \$148 \$925 \$1332 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4361 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4362 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4363 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4364 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4365 \$1333 \$265 \$265 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4366 VSS \$265 \$1333 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4367 \$1334 \$265 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4368 \$34 \$265 \$1334 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4369 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4370 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4371 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4372 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4373 \$1335 \$268 \$182 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4374 \$875 \$268 \$1335 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4375 \$1336 \$926 \$875 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4376 \$927 \$926 \$1336 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4377 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4378 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4379 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4380 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4381 \$1337 \$927 \$126 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4382 \$268 \$927 \$1337 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4383 \$1338 \$927 \$268 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4384 \$155 \$927 \$1338 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4385 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4386 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4387 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4388 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4389 \$1339 \$267 \$267 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4390 VSS \$267 \$1339 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4391 \$1340 \$267 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4392 \$35 \$267 \$1340 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4393 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4394 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4395 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4396 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4397 \$1341 \$270 \$184 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4398 \$876 \$270 \$1341 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4399 \$1342 \$928 \$876 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4400 \$929 \$928 \$1342 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4401 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4402 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4403 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4404 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4405 \$1343 \$929 \$127 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4406 \$270 \$929 \$1343 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4407 \$1344 \$929 \$270 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4408 \$162 \$929 \$1344 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4409 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4410 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4411 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4412 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4413 \$1345 \$269 \$269 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4414 VSS \$269 \$1345 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4415 \$1346 \$269 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4416 \$36 \$269 \$1346 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4417 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4418 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4419 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4420 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4421 \$1347 \$272 \$186 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4422 \$877 \$272 \$1347 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4423 \$1348 \$930 \$877 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4424 \$931 \$930 \$1348 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4425 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4426 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4427 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4428 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4429 \$1349 \$931 \$128 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4430 \$272 \$931 \$1349 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4431 \$1350 \$931 \$272 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4432 \$169 \$931 \$1350 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4433 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4434 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4435 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4436 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4437 \$1351 \$271 \$271 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4438 VSS \$271 \$1351 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4439 \$1352 \$271 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4440 \$37 \$271 \$1352 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4441 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4442 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4443 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4444 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4445 \$1353 \$274 \$188 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4446 \$878 \$274 \$1353 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4447 \$1354 \$932 \$878 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4448 \$933 \$932 \$1354 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4449 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4450 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4451 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4452 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4453 \$1355 \$933 \$129 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4454 \$274 \$933 \$1355 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4455 \$1356 \$933 \$274 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4456 \$176 \$933 \$1356 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4457 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4458 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4459 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4460 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4461 \$1357 \$273 \$273 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4462 VSS \$273 \$1357 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4463 \$1358 \$273 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4464 \$38 \$273 \$1358 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4465 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4466 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4467 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4468 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4469 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4470 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4471 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4472 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4473 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4474 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4475 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4476 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4477 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4478 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4479 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4480 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4481 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4482 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4483 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4484 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4485 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4486 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4487 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4488 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4489 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4490 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4491 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4492 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4493 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4494 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4495 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4496 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4497 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4498 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4499 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4500 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4501 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4502 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4503 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4504 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4505 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4506 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4507 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4508 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4509 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4510 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4511 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4512 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4513 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4514 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4515 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4516 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4517 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4518 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4519 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4520 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4521 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4522 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4523 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4524 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4525 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4526 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4527 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4528 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4529 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4530 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4531 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4532 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4533 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4534 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4535 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4536 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4537 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4538 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4539 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4540 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4541 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4542 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4543 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4544 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4545 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4546 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4547 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4548 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4549 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4550 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4551 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4552 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4553 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4554 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4555 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4556 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4557 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4558 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4559 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4560 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4561 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4562 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4563 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4564 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4565 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4566 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4567 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4568 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4569 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4570 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4571 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4572 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4573 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4574 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4575 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4576 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4577 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4578 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4579 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4580 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4581 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4582 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4583 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4584 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4585 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4586 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4587 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4588 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4589 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4590 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4591 \$1796 \$1769 \$1795 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4592 \$924 \$1769 \$1796 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4593 \$1798 \$1769 \$1797 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4594 \$1799 \$1769 \$1798 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4595 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4596 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4597 \$1800 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4598 \$1801 \$1769 \$1800 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4599 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4600 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4601 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4602 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4603 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4604 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4605 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4606 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4607 \$1803 \$1769 \$1802 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4608 \$926 \$1769 \$1803 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4609 \$1805 \$1769 \$1804 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4610 \$1806 \$1769 \$1805 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4611 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4612 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4613 \$1807 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4614 \$1808 \$1769 \$1807 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4615 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4616 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4617 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4618 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4619 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4620 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4621 \$1810 \$1769 \$1809 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4622 \$928 \$1769 \$1810 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4623 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4624 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4625 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4626 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4627 \$1812 \$1769 \$1811 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4628 \$1813 \$1769 \$1812 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4629 \$1814 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4630 \$1815 \$1769 \$1814 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4631 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4632 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4633 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4634 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4635 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4636 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4637 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4638 \$1966 \$1770 \$1816 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4639 \$1967 \$1770 \$1966 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4640 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4641 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4642 \$1817 \$1770 \$1816 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4643 \$1771 \$1770 \$1817 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4644 \$1969 \$1770 \$1968 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4645 \$1819 \$1770 \$1969 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4646 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4647 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4648 \$1818 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4649 \$1819 \$1770 \$1818 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4650 \$1971 \$1770 \$1970 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4651 \$1821 \$1770 \$1971 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4652 \$1820 \$1770 \$1771 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4653 \$1821 \$1770 \$1820 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4654 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4655 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4656 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4657 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4658 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4659 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4660 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4661 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4662 \$1972 \$1770 \$1822 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4663 \$1973 \$1770 \$1972 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4664 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4665 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4666 \$1823 \$1770 \$1822 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4667 \$1772 \$1770 \$1823 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4668 \$1824 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4669 \$1825 \$1770 \$1824 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4670 \$1975 \$1770 \$1974 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4671 \$1825 \$1770 \$1975 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4672 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4673 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4674 \$1977 \$1770 \$1976 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4675 \$1827 \$1770 \$1977 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4676 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4677 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4678 \$1826 \$1770 \$1772 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4679 \$1827 \$1770 \$1826 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4680 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4681 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4682 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4683 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4684 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4685 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4686 \$1829 \$1770 \$1828 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4687 \$1773 \$1770 \$1829 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4688 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4689 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4690 \$1978 \$1770 \$1828 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4691 \$1979 \$1770 \$1978 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4692 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4693 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4694 \$1981 \$1770 \$1980 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4695 \$1831 \$1770 \$1981 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4696 \$1830 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4697 \$1831 \$1770 \$1830 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4698 \$1832 \$1770 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4699 \$1833 \$1770 \$1832 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4700 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4701 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4702 \$1983 \$1770 \$1982 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4703 \$1833 \$1770 \$1983 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4704 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4705 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4706 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4707 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4708 \$1948 \$1769 \$1795 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4709 \$1949 \$1769 \$1948 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4710 \$1951 \$1769 \$1950 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4711 \$1799 \$1769 \$1951 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4712 \$1953 \$1769 \$1952 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4713 \$1801 \$1769 \$1953 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4714 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4715 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4716 \$1954 \$1769 \$1802 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4717 \$1955 \$1769 \$1954 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4718 \$1957 \$1769 \$1956 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4719 \$1806 \$1769 \$1957 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4720 \$1959 \$1769 \$1958 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4721 \$1808 \$1769 \$1959 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4722 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4723 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4724 \$1960 \$1769 \$1809 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4725 \$1961 \$1769 \$1960 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4726 \$1963 \$1769 \$1962 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4727 \$1813 \$1769 \$1963 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4728 \$1965 \$1769 \$1964 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4729 \$1815 \$1769 \$1965 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4730 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4731 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4732 \$2122 \$1769 \$2121 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4733 \$1949 \$1769 \$2122 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4734 \$2123 \$1769 \$1950 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4735 \$2124 \$1769 \$2123 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4736 \$2125 \$1769 \$1952 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4737 \$2126 \$1769 \$2125 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4738 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4739 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4740 \$2128 \$1769 \$2127 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4741 \$1955 \$1769 \$2128 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4742 \$2129 \$1769 \$1956 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4743 \$2130 \$1769 \$2129 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4744 \$2131 \$1769 \$1958 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4745 \$2132 \$1769 \$2131 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4746 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4747 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4748 \$2134 \$1769 \$2133 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4749 \$1961 \$1769 \$2134 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4750 \$2135 \$1769 \$1962 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4751 \$2136 \$1769 \$2135 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4752 \$2137 \$1769 \$1964 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4753 \$2138 \$1769 \$2137 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4754 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4755 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4756 \$2140 \$1770 \$2139 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4757 \$1967 \$1770 \$2140 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4758 \$2141 \$1770 \$1968 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4759 \$2096 \$1770 \$2141 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4760 \$2142 \$1770 \$1970 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4761 \$2143 \$1770 \$2142 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4762 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4763 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4764 \$2145 \$1770 \$2144 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4765 \$1973 \$1770 \$2145 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4766 \$2146 \$1770 \$1974 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4767 \$2097 \$1770 \$2146 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4768 \$2147 \$1770 \$1976 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4769 \$2148 \$1770 \$2147 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4770 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4771 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4772 \$2150 \$1770 \$2149 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4773 \$1979 \$1770 \$2150 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4774 \$2151 \$1770 \$1980 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4775 \$2098 \$1770 \$2151 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4776 \$2152 \$1770 \$1982 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4777 \$2153 \$1770 \$2152 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4778 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4779 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4780 \$2441 \$1769 \$2121 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4781 \$2442 \$1769 \$2441 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4782 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4783 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4784 \$2444 \$1769 \$2443 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4785 \$2126 \$1769 \$2444 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4786 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4787 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4788 \$2445 \$1769 \$2127 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4789 \$2446 \$1769 \$2445 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4790 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4791 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4792 \$2448 \$1769 \$2447 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4793 \$2132 \$1769 \$2448 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4794 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4795 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4796 \$2449 \$1769 \$2133 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4797 \$2450 \$1769 \$2449 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4798 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4799 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4800 \$2452 \$1769 \$2451 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4801 \$2138 \$1769 \$2452 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4802 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4803 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4804 \$2399 \$1770 \$2139 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4805 \$2400 \$1770 \$2399 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4806 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4807 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4808 \$2402 \$1770 \$2401 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4809 \$2143 \$1770 \$2402 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4810 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4811 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4812 \$2403 \$1770 \$2144 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4813 \$2404 \$1770 \$2403 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4814 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4815 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4816 \$2406 \$1770 \$2405 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4817 \$2148 \$1770 \$2406 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4818 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4819 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4820 \$2407 \$1770 \$2149 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4821 \$2408 \$1770 \$2407 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4822 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4823 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4824 \$2410 \$1770 \$2409 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4825 \$2153 \$1770 \$2410 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4826 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4827 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4828 \$2696 \$1769 \$874 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4829 \$1797 \$1769 \$2696 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4830 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4831 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4832 \$2697 \$1769 \$2124 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4833 \$2698 \$1769 \$2697 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4834 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4835 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4836 \$2699 \$1769 \$875 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4837 \$1804 \$1769 \$2699 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4838 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4839 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4840 \$2700 \$1769 \$2130 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4841 \$2701 \$1769 \$2700 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4842 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4843 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4844 \$2702 \$1769 \$876 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4845 \$1811 \$1769 \$2702 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4846 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4847 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4848 \$2703 \$1769 \$2136 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4849 \$2704 \$1769 \$2703 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4850 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4851 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4852 \$2705 \$1770 \$5667 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4853 \$2706 \$1770 \$2705 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4854 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4855 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4856 \$2708 \$1770 \$2707 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4857 \$2096 \$1770 \$2708 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4858 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4859 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4860 \$2709 \$1770 \$5668 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4861 \$2710 \$1770 \$2709 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4862 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4863 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4864 \$2712 \$1770 \$2711 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4865 \$2097 \$1770 \$2712 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4866 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4867 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4868 \$2713 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4869 \$2714 \$1770 \$2713 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4870 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4871 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4872 \$2716 \$1770 \$2715 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4873 \$2098 \$1770 \$2716 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4874 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4875 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4876 \$2938 \$1769 \$2937 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4877 \$2442 \$1769 \$2938 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4878 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4879 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4880 \$2939 \$1769 \$2443 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4881 \$2940 \$1769 \$2939 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4882 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4883 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4884 \$2942 \$1769 \$2941 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4885 \$2446 \$1769 \$2942 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4886 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4887 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4888 \$2943 \$1769 \$2447 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4889 \$2944 \$1769 \$2943 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4890 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4891 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4892 \$2946 \$1769 \$2945 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4893 \$2450 \$1769 \$2946 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4894 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4895 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4896 \$2947 \$1769 \$2451 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4897 \$2948 \$1769 \$2947 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4898 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4899 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4900 \$2950 \$1770 \$2949 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4901 \$2400 \$1770 \$2950 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4902 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4903 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4904 \$2951 \$1770 \$2401 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4905 \$2952 \$1770 \$2951 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4906 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4907 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4908 \$2954 \$1770 \$2953 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4909 \$2404 \$1770 \$2954 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4910 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4911 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4912 \$2955 \$1770 \$2405 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4913 \$2956 \$1770 \$2955 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4914 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4915 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4916 \$2958 \$1770 \$2957 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4917 \$2408 \$1770 \$2958 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4918 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4919 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4920 \$2959 \$1770 \$2409 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4921 \$2960 \$1770 \$2959 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4922 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4923 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4924 \$3207 \$1769 \$2937 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4925 \$3208 \$1769 \$3207 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4926 \$3210 \$1769 \$3209 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4927 \$2698 \$1769 \$3210 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4928 \$3212 \$1769 \$3211 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4929 \$2940 \$1769 \$3212 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4930 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4931 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4932 \$3213 \$1769 \$2941 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4933 \$3214 \$1769 \$3213 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4934 \$3216 \$1769 \$3215 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4935 \$2701 \$1769 \$3216 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4936 \$3218 \$1769 \$3217 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4937 \$2944 \$1769 \$3218 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4938 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4939 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4940 \$3219 \$1769 \$2945 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4941 \$3220 \$1769 \$3219 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4942 \$3222 \$1769 \$3221 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4943 \$2704 \$1769 \$3222 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4944 \$3224 \$1769 \$3223 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4945 \$2948 \$1769 \$3224 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4946 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4947 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4948 \$3225 \$1770 \$2949 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4949 \$3226 \$1770 \$3225 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4950 \$3228 \$1770 \$3227 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4951 \$2707 \$1770 \$3228 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4952 \$3230 \$1770 \$3229 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4953 \$2952 \$1770 \$3230 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4954 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4955 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4956 \$3231 \$1770 \$2953 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4957 \$3232 \$1770 \$3231 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4958 \$3234 \$1770 \$3233 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4959 \$2711 \$1770 \$3234 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4960 \$3236 \$1770 \$3235 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4961 \$2956 \$1770 \$3236 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4962 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4963 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4964 \$3237 \$1770 \$2957 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4965 \$3238 \$1770 \$3237 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4966 \$3240 \$1770 \$3239 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4967 \$2715 \$1770 \$3240 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4968 \$3242 \$1770 \$3241 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4969 \$2960 \$1770 \$3242 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4970 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4971 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4972 \$3506 \$1769 \$3505 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4973 \$3208 \$1769 \$3506 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4974 \$3507 \$1769 \$3209 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4975 \$3508 \$1769 \$3507 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4976 \$3509 \$1769 \$3211 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4977 \$3510 \$1769 \$3509 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4978 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4979 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4980 \$3512 \$1769 \$3511 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4981 \$3214 \$1769 \$3512 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4982 \$3513 \$1769 \$3215 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4983 \$3514 \$1769 \$3513 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4984 \$3515 \$1769 \$3217 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4985 \$3516 \$1769 \$3515 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4986 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4987 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4988 \$3518 \$1769 \$3517 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4989 \$3220 \$1769 \$3518 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4990 \$3519 \$1769 \$3221 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4991 \$3520 \$1769 \$3519 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4992 \$3521 \$1769 \$3223 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4993 \$3522 \$1769 \$3521 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4994 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4995 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4996 \$3524 \$1770 \$3523 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4997 \$3226 \$1770 \$3524 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4998 \$3525 \$1770 \$3227 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4999 \$3526 \$1770 \$3525 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5000 \$3527 \$1770 \$3229 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5001 \$3528 \$1770 \$3527 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5002 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5003 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5004 \$3530 \$1770 \$3529 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5005 \$3232 \$1770 \$3530 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5006 \$3531 \$1770 \$3233 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5007 \$3532 \$1770 \$3531 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5008 \$3533 \$1770 \$3235 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5009 \$3534 \$1770 \$3533 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5010 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5011 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5012 \$3536 \$1770 \$3535 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5013 \$3238 \$1770 \$3536 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5014 \$3537 \$1770 \$3239 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5015 \$3538 \$1770 \$3537 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5016 \$3539 \$1770 \$3241 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5017 \$3540 \$1770 \$3539 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5018 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5019 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5020 \$3654 \$1769 \$3505 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5021 \$3655 \$1769 \$3654 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5022 \$3656 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5023 \$3508 \$1769 \$3656 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5024 \$3657 \$1769 \$3655 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5025 \$3510 \$1769 \$3657 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5026 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5027 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5028 \$3658 \$1769 \$3511 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5029 \$3659 \$1769 \$3658 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5030 \$3660 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5031 \$3514 \$1769 \$3660 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5032 \$3661 \$1769 \$3659 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5033 \$3516 \$1769 \$3661 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5034 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5035 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5036 \$3662 \$1769 \$3517 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5037 \$3663 \$1769 \$3662 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5038 \$3664 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5039 \$3520 \$1769 \$3664 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5040 \$3665 \$1769 \$3663 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5041 \$3522 \$1769 \$3665 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5042 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5043 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5044 \$3666 \$1770 \$3523 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5045 \$3667 \$1770 \$3666 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5046 \$3668 \$1770 \$2706 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5047 \$3526 \$1770 \$3668 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5048 \$3669 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5049 \$3528 \$1770 \$3669 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5050 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5051 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5052 \$3670 \$1770 \$3529 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5053 \$3671 \$1770 \$3670 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5054 \$3672 \$1770 \$2710 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5055 \$3532 \$1770 \$3672 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5056 \$3673 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5057 \$3534 \$1770 \$3673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5058 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5059 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5060 \$3674 \$1770 \$3535 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5061 IBNOUT \$1770 \$3674 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5062 \$3676 \$1770 \$2714 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5063 \$3538 \$1770 \$3676 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5064 \$3677 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5065 \$3540 \$1770 \$3677 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5066 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5067 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5068 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5069 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5070 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5071 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5072 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5073 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5074 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5075 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5076 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5077 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5078 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5079 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5080 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5081 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5082 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5083 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5084 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5085 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5086 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5087 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5088 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5089 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5090 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5091 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5092 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5093 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5094 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5095 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5096 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5097 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5098 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5099 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5100 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5101 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5102 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5103 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5104 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5105 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5106 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5107 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5108 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5109 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5110 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5111 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5112 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5113 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5114 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5115 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5116 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5117 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5118 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5119 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5120 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5121 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5122 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5123 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5124 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5125 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5126 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5127 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5128 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5129 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5130 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5131 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5132 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5133 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5134 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5135 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5136 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5137 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5138 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5139 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5140 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5141 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5142 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5143 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5144 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5145 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5146 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5147 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5148 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5149 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5150 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5151 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5152 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5153 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5154 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5155 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5156 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5157 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5158 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5159 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5160 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5161 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5162 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5163 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5164 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5165 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5166 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5167 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5168 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5169 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5170 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5171 \$3778 I1N I1N VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5172 VSS I1N \$3778 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5173 \$3866 I1N \$1581 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5174 VSS I1N \$3866 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5175 \$3779 I1N VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5176 \$1582 I1N \$3779 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5177 \$3867 I1N VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5178 \$4700 I1N \$3867 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5179 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5180 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5181 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5182 \$4034 \$1769 \$4033 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5183 \$930 \$1769 \$4034 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5184 \$4036 \$1769 \$4035 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5185 \$4037 \$1769 \$4036 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5186 \$4038 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5187 \$4039 \$1769 \$4038 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5188 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5189 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5190 \$4041 \$1769 \$4040 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5191 \$932 \$1769 \$4041 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5192 \$4043 \$1769 \$4042 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5193 \$4044 \$1769 \$4043 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5194 \$4045 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5195 \$4046 \$1769 \$4045 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5196 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5197 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5198 \$4048 \$1769 \$4047 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5199 VSS \$1769 \$4048 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5200 \$4050 \$1769 \$4049 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5201 \$4051 \$1769 \$4050 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5202 \$4052 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5203 \$4053 \$1769 \$4052 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5204 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5205 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5206 \$4003 \$1770 \$4002 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5207 \$3946 \$1770 \$4003 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5208 \$4004 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5209 \$4005 \$1770 \$4004 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5210 \$4006 \$1770 \$3946 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5211 \$4007 \$1770 \$4006 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5212 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5213 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5214 \$4009 \$1770 \$4008 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5215 \$3947 \$1770 \$4009 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5216 \$4010 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5217 \$4011 \$1770 \$4010 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5218 \$4012 \$1770 \$3947 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5219 \$4013 \$1770 \$4012 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5220 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5221 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5222 \$4015 \$1770 \$4014 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5223 \$3948 \$1770 \$4015 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5224 \$4016 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5225 \$4017 \$1770 \$4016 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5226 \$4018 \$1770 \$3948 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5227 \$4019 \$1770 \$4018 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5228 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5229 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5230 \$3949 I1N \$1581 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5231 VSS I1N \$3949 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5232 \$3950 I1N VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5233 \$4700 I1N \$3950 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5234 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5235 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5236 \$4183 \$1769 \$4033 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5237 \$4184 \$1769 \$4183 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5238 \$4186 \$1769 \$4185 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5239 \$4037 \$1769 \$4186 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5240 \$4188 \$1769 \$4187 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5241 \$4039 \$1769 \$4188 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5242 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5243 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5244 \$4189 \$1769 \$4040 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5245 \$4190 \$1769 \$4189 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5246 \$4192 \$1769 \$4191 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5247 \$4044 \$1769 \$4192 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5248 \$4194 \$1769 \$4193 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5249 \$4046 \$1769 \$4194 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5250 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5251 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5252 \$4195 \$1769 \$4047 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5253 \$4196 \$1769 \$4195 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5254 \$4198 \$1769 \$4197 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5255 \$4051 \$1769 \$4198 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5256 \$4200 \$1769 \$4199 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5257 \$4053 \$1769 \$4200 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5258 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5259 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5260 \$4201 \$1770 \$4002 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5261 \$4202 \$1770 \$4201 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5262 \$4204 \$1770 \$4203 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5263 \$4005 \$1770 \$4204 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5264 \$4206 \$1770 \$4205 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5265 \$4007 \$1770 \$4206 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5266 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5267 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5268 \$4207 \$1770 \$4008 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5269 \$4208 \$1770 \$4207 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5270 \$4210 \$1770 \$4209 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5271 \$4011 \$1770 \$4210 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5272 \$4212 \$1770 \$4211 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5273 \$4013 \$1770 \$4212 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5274 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5275 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5276 \$4213 \$1770 \$4014 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5277 \$4214 \$1770 \$4213 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5278 \$4216 \$1770 \$4215 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5279 \$4017 \$1770 \$4216 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5280 \$4218 \$1770 \$4217 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5281 \$4019 \$1770 \$4218 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5282 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5283 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5284 \$4098 I1N \$1582 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5285 VSS I1N \$4098 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5286 \$4099 I1N VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5287 I1N I1N \$4099 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5288 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5289 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5290 \$4343 \$1769 \$4342 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5291 \$4184 \$1769 \$4343 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5292 \$4344 \$1769 \$4185 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5293 \$4345 \$1769 \$4344 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5294 \$4346 \$1769 \$4187 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5295 \$4347 \$1769 \$4346 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5296 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5297 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5298 \$4349 \$1769 \$4348 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5299 \$4190 \$1769 \$4349 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5300 \$4350 \$1769 \$4191 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5301 \$4351 \$1769 \$4350 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5302 \$4352 \$1769 \$4193 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5303 \$4353 \$1769 \$4352 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5304 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5305 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5306 \$4355 \$1769 \$4354 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5307 \$4196 \$1769 \$4355 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5308 \$4356 \$1769 \$4197 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5309 \$4357 \$1769 \$4356 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5310 \$4358 \$1769 \$4199 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5311 \$4359 \$1769 \$4358 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5312 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5313 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5314 \$4361 \$1770 \$4360 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5315 \$4202 \$1770 \$4361 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5316 \$4362 \$1770 \$4203 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5317 \$4257 \$1770 \$4362 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5318 \$4363 \$1770 \$4205 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5319 \$4364 \$1770 \$4363 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5320 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5321 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5322 \$4366 \$1770 \$4365 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5323 \$4208 \$1770 \$4366 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5324 \$4367 \$1770 \$4209 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5325 \$4258 \$1770 \$4367 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5326 \$4368 \$1770 \$4211 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5327 \$4369 \$1770 \$4368 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5328 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5329 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5330 \$4371 \$1770 \$4370 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5331 \$4214 \$1770 \$4371 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5332 \$4372 \$1770 \$4215 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5333 \$4259 \$1770 \$4372 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5334 \$4373 \$1770 \$4217 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5335 \$4374 \$1770 \$4373 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5336 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5337 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5338 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5339 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5340 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5341 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5342 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5343 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5344 \$4515 \$1769 \$4342 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5345 \$4516 \$1769 \$4515 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5346 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5347 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5348 \$4518 \$1769 \$4517 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5349 \$4347 \$1769 \$4518 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5350 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5351 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5352 \$4519 \$1769 \$4348 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5353 \$4520 \$1769 \$4519 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5354 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5355 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5356 \$4522 \$1769 \$4521 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5357 \$4353 \$1769 \$4522 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5358 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5359 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5360 \$4523 \$1769 \$4354 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5361 \$4524 \$1769 \$4523 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5362 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5363 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5364 \$4526 \$1769 \$4525 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5365 \$4359 \$1769 \$4526 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5366 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5367 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5368 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5369 \$4688 \$1770 \$5664 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5370 \$4689 \$1770 \$4688 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5371 \$4527 \$1770 \$4360 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5372 \$4528 \$1770 \$4527 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5373 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5374 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5375 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5376 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5377 \$4530 \$1770 \$4529 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5378 \$4364 \$1770 \$4530 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5379 \$4690 \$1770 \$4697 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5380 \$4257 \$1770 \$4690 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5381 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5382 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5383 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5384 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5385 \$4691 \$1770 \$5665 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5386 \$4692 \$1770 \$4691 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5387 \$4531 \$1770 \$4365 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5388 \$4532 \$1770 \$4531 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5389 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5390 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5391 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5392 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5393 \$4534 \$1770 \$4533 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5394 \$4369 \$1770 \$4534 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5395 \$4693 \$1770 \$4698 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5396 \$4258 \$1770 \$4693 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5397 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5398 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5399 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5400 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5401 \$4694 \$1770 \$5666 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5402 \$4695 \$1770 \$4694 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5403 \$4535 \$1770 \$4370 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5404 \$4536 \$1770 \$4535 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5405 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5406 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5407 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5408 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5409 \$4538 \$1770 \$4537 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5410 \$4374 \$1770 \$4538 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5411 \$4696 \$1770 \$4699 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5412 \$4259 \$1770 \$4696 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5413 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5414 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5415 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5416 \$4679 \$1769 \$877 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5417 \$4035 \$1769 \$4679 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5418 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5419 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5420 \$4680 \$1769 \$4345 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5421 \$4681 \$1769 \$4680 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5422 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5423 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5424 \$4682 \$1769 \$878 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5425 \$4042 \$1769 \$4682 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5426 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5427 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5428 \$4683 \$1769 \$4351 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5429 \$4684 \$1769 \$4683 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5430 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5431 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5432 \$4685 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5433 \$4049 \$1769 \$4685 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5434 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5435 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5436 \$4686 \$1769 \$4357 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5437 \$4687 \$1769 \$4686 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5438 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5439 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5440 \$4839 \$1769 \$4838 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5441 \$4516 \$1769 \$4839 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5442 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5443 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5444 \$4840 \$1769 \$4517 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5445 \$4841 \$1769 \$4840 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5446 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5447 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5448 \$4843 \$1769 \$4842 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5449 \$4520 \$1769 \$4843 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5450 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5451 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5452 \$4844 \$1769 \$4521 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5453 \$4845 \$1769 \$4844 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5454 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5455 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5456 \$4847 \$1769 \$4846 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5457 \$4524 \$1769 \$4847 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5458 VSS \$1769 \$1769 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5459 \$1769 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5460 \$4848 \$1769 \$4525 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5461 \$4849 \$1769 \$4848 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5462 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5463 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5464 \$4851 \$1770 \$4850 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5465 \$4528 \$1770 \$4851 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5466 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5467 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5468 \$4852 \$1770 \$4529 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5469 \$4853 \$1770 \$4852 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5470 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5471 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5472 \$4855 \$1770 \$4854 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5473 \$4532 \$1770 \$4855 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5474 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5475 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5476 \$4856 \$1770 \$4533 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5477 \$4857 \$1770 \$4856 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5478 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5479 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5480 \$4859 \$1770 \$4858 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5481 \$4536 \$1770 \$4859 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5482 VSS \$1770 \$1770 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5483 \$1770 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5484 \$4860 \$1770 \$4537 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5485 \$4861 \$1770 \$4860 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5486 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5487 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5488 \$5040 \$1769 \$4838 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5489 \$5041 \$1769 \$5040 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5490 \$5043 \$1769 \$5042 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5491 \$4681 \$1769 \$5043 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5492 \$5045 \$1769 \$5044 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5493 \$4841 \$1769 \$5045 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5494 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5495 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5496 \$5046 \$1769 \$4842 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5497 \$5047 \$1769 \$5046 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5498 \$5049 \$1769 \$5048 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5499 \$4684 \$1769 \$5049 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5500 \$5051 \$1769 \$5050 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5501 \$4845 \$1769 \$5051 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5502 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5503 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5504 \$5052 \$1769 \$4846 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5505 \$5053 \$1769 \$5052 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5506 \$5055 \$1769 \$5054 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5507 \$4687 \$1769 \$5055 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5508 \$5057 \$1769 \$5056 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5509 \$4849 \$1769 \$5057 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5510 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5511 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5512 \$5011 \$1770 \$4850 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5513 \$5012 \$1770 \$5011 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5514 \$5014 \$1770 \$5013 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5515 \$4697 \$1770 \$5014 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5516 \$5016 \$1770 \$5015 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5517 \$4853 \$1770 \$5016 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5518 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5519 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5520 \$5017 \$1770 \$4854 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5521 \$5018 \$1770 \$5017 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5522 \$5020 \$1770 \$5019 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5523 \$4698 \$1770 \$5020 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5524 \$5022 \$1770 \$5021 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5525 \$4857 \$1770 \$5022 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5526 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5527 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5528 \$5023 \$1770 \$4858 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5529 \$5024 \$1770 \$5023 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5530 \$5026 \$1770 \$5025 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5531 \$4699 \$1770 \$5026 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5532 \$5028 \$1770 \$5027 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5533 \$4861 \$1770 \$5028 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5534 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5535 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5536 \$5187 \$1769 \$5186 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5537 \$5041 \$1769 \$5187 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5538 \$5188 \$1769 \$5042 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5539 \$5189 \$1769 \$5188 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5540 \$5190 \$1769 \$5044 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5541 \$5191 \$1769 \$5190 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5542 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5543 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5544 \$5193 \$1769 \$5192 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5545 \$5047 \$1769 \$5193 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5546 \$5194 \$1769 \$5048 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5547 \$5195 \$1769 \$5194 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5548 \$5196 \$1769 \$5050 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5549 \$5197 \$1769 \$5196 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5550 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5551 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5552 \$5199 \$1769 \$5198 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5553 \$5053 \$1769 \$5199 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5554 \$5200 \$1769 \$5054 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5555 \$5201 \$1769 \$5200 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5556 \$5202 \$1769 \$5056 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5557 \$5203 \$1769 \$5202 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5558 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5559 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5560 \$5205 \$1770 \$5204 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5561 \$5012 \$1770 \$5205 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5562 \$5206 \$1770 \$5013 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5563 \$5207 \$1770 \$5206 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5564 \$5208 \$1770 \$5015 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5565 \$5209 \$1770 \$5208 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5566 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5567 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5568 \$5211 \$1770 \$5210 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5569 \$5018 \$1770 \$5211 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5570 \$5212 \$1770 \$5019 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5571 \$5213 \$1770 \$5212 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5572 \$5214 \$1770 \$5021 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5573 \$5215 \$1770 \$5214 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5574 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5575 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5576 \$5217 \$1770 \$5216 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5577 \$5024 \$1770 \$5217 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5578 \$5218 \$1770 \$5025 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5579 \$5219 \$1770 \$5218 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5580 \$5220 \$1770 \$5027 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5581 \$5221 \$1770 \$5220 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5582 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5583 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5584 \$5327 \$1769 \$5186 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5585 \$5328 \$1769 \$5327 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5586 \$5329 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5587 \$5189 \$1769 \$5329 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5588 \$5330 \$1769 \$5328 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5589 \$5191 \$1769 \$5330 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5590 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5591 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5592 \$5331 \$1769 \$5192 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5593 \$5332 \$1769 \$5331 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5594 \$5333 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5595 \$5195 \$1769 \$5333 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5596 \$5334 \$1769 \$5332 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5597 \$5197 \$1769 \$5334 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5598 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5599 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5600 \$5335 \$1769 \$5198 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5601 \$5336 \$1769 \$5335 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5602 \$5337 \$1769 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5603 \$5201 \$1769 \$5337 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5604 \$5338 \$1769 \$5336 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5605 \$5203 \$1769 \$5338 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5606 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5607 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5608 \$5339 \$1770 \$5204 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5609 \$5340 \$1770 \$5339 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5610 \$5341 \$1770 \$4689 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5611 \$5207 \$1770 \$5341 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5612 \$5342 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5613 \$5209 \$1770 \$5342 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5614 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5615 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5616 \$5343 \$1770 \$5210 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5617 \$5344 \$1770 \$5343 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5618 \$5345 \$1770 \$4692 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5619 \$5213 \$1770 \$5345 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5620 \$5346 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5621 \$5215 \$1770 \$5346 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5622 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5623 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5624 \$5347 \$1770 \$5216 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5625 \$5348 \$1770 \$5347 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5626 \$5349 \$1770 \$4695 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5627 \$5219 \$1770 \$5349 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5628 \$5350 \$1770 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5629 \$5221 \$1770 \$5350 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5630 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5631 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5632 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5633 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5634 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5635 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5636 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5637 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5638 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5639 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5640 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5641 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5642 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5643 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5644 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5645 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5646 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5647 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5648 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5649 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5650 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5651 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5652 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5653 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5654 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5655 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5656 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5657 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5658 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5659 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5660 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5661 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5662 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5663 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5664 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5665 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5666 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5667 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5668 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5669 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5670 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5671 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5672 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5673 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5674 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5675 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5676 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5677 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5678 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5679 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5680 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5681 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5682 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5683 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5684 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5685 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5686 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5687 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5688 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5689 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5690 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5691 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5692 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5693 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5694 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5695 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5696 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5697 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5698 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5699 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5700 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5701 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5702 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5703 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5704 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5705 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5706 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5707 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5708 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5709 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5710 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5711 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5712 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5713 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5714 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5715 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5716 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5717 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5718 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5719 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5720 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5721 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5722 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5723 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5724 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5725 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5726 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5727 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5728 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5729 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5730 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5731 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5732 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5733 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5734 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5735 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5736 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5737 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5738 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5739 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5740 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5741 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5742 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5743 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5744 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5745 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5746 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5747 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5748 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5749 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5750 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5751 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5752 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5753 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5754 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5755 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5756 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5757 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5758 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5759 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5760 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5761 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5762 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5763 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5764 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5765 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5766 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5767 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5768 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5769 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5770 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5771 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5772 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5773 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5774 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5775 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5776 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5777 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5778 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5779 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5780 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5781 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5782 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5783 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5784 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5785 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5786 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5787 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5788 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5789 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5790 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5791 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5792 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5793 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5794 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5795 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5796 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5797 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5798 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5799 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5800 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5801 \$5690 \$5789 \$5689 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5802 \$5664 \$5789 \$5690 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5803 \$5691 \$5340 \$5664 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5804 \$5588 \$5340 \$5691 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5805 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5806 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5807 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5808 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5809 \$5693 \$5588 \$5692 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5810 \$5789 \$5588 \$5693 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5811 \$5694 \$5588 \$5789 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5812 \$5799 \$5588 \$5694 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5813 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5814 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5815 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5816 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5817 \$5695 \$5790 \$5790 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5818 VSS \$5790 \$5695 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5819 \$5696 \$5790 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5820 \$6468 \$5790 \$5696 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5821 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5822 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5823 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5824 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5825 \$5698 \$5791 \$5697 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5826 \$5665 \$5791 \$5698 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5827 \$5699 \$5344 \$5665 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5828 \$5589 \$5344 \$5699 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5829 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5830 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5831 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5832 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5833 \$5701 \$5589 \$5700 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5834 \$5791 \$5589 \$5701 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5835 \$5702 \$5589 \$5791 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5836 \$5800 \$5589 \$5702 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5837 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5838 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5839 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5840 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5841 \$5703 \$5792 \$5792 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5842 VSS \$5792 \$5703 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5843 \$5704 \$5792 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5844 \$6469 \$5792 \$5704 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5845 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5846 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5847 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5848 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5849 \$5706 \$5793 \$5705 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5850 \$5666 \$5793 \$5706 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5851 \$5707 \$5348 \$5666 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5852 \$5590 \$5348 \$5707 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5853 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5854 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5855 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5856 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5857 \$5709 \$5590 \$5708 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5858 \$5793 \$5590 \$5709 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5859 \$5710 \$5590 \$5793 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5860 \$5801 \$5590 \$5710 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5861 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5862 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5863 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5864 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5865 \$5711 \$5794 \$5794 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5866 VSS \$5794 \$5711 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5867 \$5712 \$5794 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5868 \$6470 \$5794 \$5712 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5869 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5870 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5871 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5872 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5873 \$5714 \$5795 \$5713 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5874 \$5667 \$5795 \$5714 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5875 \$5715 \$3667 \$5667 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5876 \$5591 \$3667 \$5715 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5877 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5878 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5879 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5880 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5881 \$5717 \$5591 \$5716 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5882 \$5795 \$5591 \$5717 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5883 \$5718 \$5591 \$5795 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5884 \$5802 \$5591 \$5718 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5885 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5886 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5887 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5888 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5889 \$5719 \$5796 \$5796 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5890 VSS \$5796 \$5719 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5891 \$5720 \$5796 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5892 \$6471 \$5796 \$5720 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5893 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5894 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5895 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5896 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5897 \$5722 \$5797 \$5721 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5898 \$5668 \$5797 \$5722 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5899 \$5723 \$3671 \$5668 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5900 \$5592 \$3671 \$5723 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5901 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5902 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5903 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5904 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5905 \$5725 \$5592 \$5724 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5906 \$5797 \$5592 \$5725 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5907 \$5726 \$5592 \$5797 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5908 \$5803 \$5592 \$5726 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5909 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5910 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5911 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5912 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5913 \$5727 \$5798 \$5798 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5914 VSS \$5798 \$5727 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5915 \$5728 \$5798 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5916 \$6472 \$5798 \$5728 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5917 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5918 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5919 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5920 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5921 \$5859 \$5340 \$5588 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5922 \$5664 \$5340 \$5859 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5923 \$5860 \$5789 \$5664 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5924 \$5689 \$5789 \$5860 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5925 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5926 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5927 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5928 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5929 \$5861 \$5588 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5930 \$5340 \$5588 \$5861 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5931 \$5862 \$5588 \$5340 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5932 VDD \$5588 \$5862 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5933 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5934 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5935 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5936 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5937 \$5863 \$5790 \$6468 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5938 VSS \$5790 \$5863 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5939 \$5864 \$5790 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5940 \$5790 \$5790 \$5864 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5941 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5942 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5943 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5944 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5945 \$5865 \$5344 \$5589 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5946 \$5665 \$5344 \$5865 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5947 \$5866 \$5791 \$5665 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5948 \$5697 \$5791 \$5866 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5949 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5950 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5951 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5952 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5953 \$5867 \$5589 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5954 \$5344 \$5589 \$5867 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5955 \$5868 \$5589 \$5344 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5956 VDD \$5589 \$5868 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5957 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5958 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5959 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5960 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5961 \$5869 \$5792 \$6469 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5962 VSS \$5792 \$5869 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5963 \$5870 \$5792 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5964 \$5792 \$5792 \$5870 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5965 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5966 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5967 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5968 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5969 \$5871 \$5348 \$5590 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5970 \$5666 \$5348 \$5871 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5971 \$5872 \$5793 \$5666 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5972 \$5705 \$5793 \$5872 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5973 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5974 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5975 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5976 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5977 \$5873 \$5590 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5978 \$5348 \$5590 \$5873 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5979 \$5874 \$5590 \$5348 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5980 VDD \$5590 \$5874 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5981 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5982 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5983 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5984 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5985 \$5875 \$5794 \$6470 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5986 VSS \$5794 \$5875 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5987 \$5876 \$5794 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5988 \$5794 \$5794 \$5876 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5989 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5990 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5991 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5992 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5993 \$5877 \$3667 \$5591 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5994 \$5667 \$3667 \$5877 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5995 \$5878 \$5795 \$5667 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5996 \$5713 \$5795 \$5878 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5997 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5998 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5999 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6000 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6001 \$5879 \$5591 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6002 \$3667 \$5591 \$5879 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6003 \$5880 \$5591 \$3667 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6004 VDD \$5591 \$5880 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6005 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6006 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6007 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6008 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6009 \$5881 \$5796 \$6471 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6010 VSS \$5796 \$5881 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6011 \$5882 \$5796 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6012 \$5796 \$5796 \$5882 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6013 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6014 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6015 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6016 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6017 \$5883 \$3671 \$5592 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6018 \$5668 \$3671 \$5883 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6019 \$5884 \$5797 \$5668 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6020 \$5721 \$5797 \$5884 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6021 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6022 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6023 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6024 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6025 \$5885 \$5592 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6026 \$3671 \$5592 \$5885 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6027 \$5886 \$5592 \$3671 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6028 VDD \$5592 \$5886 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6029 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6030 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6031 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6032 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6033 \$5887 \$5798 \$6472 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6034 VSS \$5798 \$5887 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6035 \$5888 \$5798 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6036 \$5798 \$5798 \$5888 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6037 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6038 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6039 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6040 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6041 \$5994 \$5789 \$5689 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6042 \$5664 \$5789 \$5994 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6043 \$5995 \$5340 \$5664 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6044 \$5588 \$5340 \$5995 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6045 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6046 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6047 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6048 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6049 \$5996 \$5588 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6050 \$5340 \$5588 \$5996 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6051 \$5997 \$5588 \$5340 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6052 VDD \$5588 \$5997 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6053 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6054 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6055 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6056 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6057 \$5998 \$5790 \$5790 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6058 VSS \$5790 \$5998 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6059 \$5999 \$5790 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6060 \$6468 \$5790 \$5999 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6061 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6062 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6063 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6064 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6065 \$6000 \$5791 \$5697 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6066 \$5665 \$5791 \$6000 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6067 \$6001 \$5344 \$5665 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6068 \$5589 \$5344 \$6001 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6069 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6070 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6071 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6072 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6073 \$6002 \$5589 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6074 \$5344 \$5589 \$6002 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6075 \$6003 \$5589 \$5344 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6076 VDD \$5589 \$6003 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6077 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6078 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6079 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6080 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6081 \$6004 \$5792 \$5792 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6082 VSS \$5792 \$6004 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6083 \$6005 \$5792 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6084 \$6469 \$5792 \$6005 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6085 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6086 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6087 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6088 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6089 \$6006 \$5793 \$5705 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6090 \$5666 \$5793 \$6006 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6091 \$6007 \$5348 \$5666 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6092 \$5590 \$5348 \$6007 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6093 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6094 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6095 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6096 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6097 \$6008 \$5590 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6098 \$5348 \$5590 \$6008 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6099 \$6009 \$5590 \$5348 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6100 VDD \$5590 \$6009 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6101 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6102 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6103 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6104 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6105 \$6010 \$5794 \$5794 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6106 VSS \$5794 \$6010 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6107 \$6011 \$5794 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6108 \$6470 \$5794 \$6011 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6109 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6110 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6111 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6112 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6113 \$6012 \$5795 \$5713 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6114 \$5667 \$5795 \$6012 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6115 \$6013 \$3667 \$5667 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6116 \$5591 \$3667 \$6013 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6117 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6118 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6119 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6120 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6121 \$6014 \$5591 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6122 \$3667 \$5591 \$6014 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6123 \$6015 \$5591 \$3667 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6124 VDD \$5591 \$6015 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6125 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6126 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6127 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6128 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6129 \$6016 \$5796 \$5796 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6130 VSS \$5796 \$6016 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6131 \$6017 \$5796 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6132 \$6471 \$5796 \$6017 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6133 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6134 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6135 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6136 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6137 \$6018 \$5797 \$5721 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6138 \$5668 \$5797 \$6018 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6139 \$6019 \$3671 \$5668 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6140 \$5592 \$3671 \$6019 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6141 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6142 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6143 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6144 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6145 \$6020 \$5592 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6146 \$3671 \$5592 \$6020 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6147 \$6021 \$5592 \$3671 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6148 VDD \$5592 \$6021 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6149 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6150 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6151 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6152 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6153 \$6022 \$5798 \$5798 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6154 VSS \$5798 \$6022 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6155 \$6023 \$5798 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6156 \$6472 \$5798 \$6023 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6157 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6158 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6159 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6160 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6161 \$6139 \$5340 \$5588 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6162 \$5664 \$5340 \$6139 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6163 \$6140 \$5789 \$5664 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6164 \$5689 \$5789 \$6140 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6165 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6166 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6167 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6168 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6169 \$6141 \$5588 \$5799 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6170 \$5789 \$5588 \$6141 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6171 \$6142 \$5588 \$5789 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6172 \$5692 \$5588 \$6142 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6173 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6174 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6175 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6176 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6177 \$6143 \$5790 \$6468 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6178 VSS \$5790 \$6143 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6179 \$6144 \$5790 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6180 \$5790 \$5790 \$6144 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6181 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6182 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6183 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6184 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6185 \$6145 \$5344 \$5589 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6186 \$5665 \$5344 \$6145 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6187 \$6146 \$5791 \$5665 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6188 \$5697 \$5791 \$6146 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6189 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6190 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6191 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6192 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6193 \$6147 \$5589 \$5800 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6194 \$5791 \$5589 \$6147 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6195 \$6148 \$5589 \$5791 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6196 \$5700 \$5589 \$6148 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6197 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6198 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6199 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6200 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6201 \$6149 \$5792 \$6469 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6202 VSS \$5792 \$6149 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6203 \$6150 \$5792 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6204 \$5792 \$5792 \$6150 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6205 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6206 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6207 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6208 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6209 \$6151 \$5348 \$5590 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6210 \$5666 \$5348 \$6151 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6211 \$6152 \$5793 \$5666 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6212 \$5705 \$5793 \$6152 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6213 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6214 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6215 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6216 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6217 \$6153 \$5590 \$5801 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6218 \$5793 \$5590 \$6153 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6219 \$6154 \$5590 \$5793 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6220 \$5708 \$5590 \$6154 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6221 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6222 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6223 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6224 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6225 \$6155 \$5794 \$6470 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6226 VSS \$5794 \$6155 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6227 \$6156 \$5794 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6228 \$5794 \$5794 \$6156 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6229 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6230 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6231 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6232 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6233 \$6157 \$3667 \$5591 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6234 \$5667 \$3667 \$6157 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6235 \$6158 \$5795 \$5667 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6236 \$5713 \$5795 \$6158 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6237 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6238 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6239 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6240 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6241 \$6159 \$5591 \$5802 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6242 \$5795 \$5591 \$6159 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6243 \$6160 \$5591 \$5795 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6244 \$5716 \$5591 \$6160 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6245 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6246 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6247 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6248 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6249 \$6161 \$5796 \$6471 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6250 VSS \$5796 \$6161 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6251 \$6162 \$5796 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6252 \$5796 \$5796 \$6162 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6253 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6254 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6255 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6256 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6257 \$6163 \$3671 \$5592 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6258 \$5668 \$3671 \$6163 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6259 \$6164 \$5797 \$5668 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6260 \$5721 \$5797 \$6164 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6261 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6262 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6263 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6264 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6265 \$6165 \$5592 \$5803 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6266 \$5797 \$5592 \$6165 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6267 \$6166 \$5592 \$5797 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6268 \$5724 \$5592 \$6166 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6269 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6270 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6271 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6272 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6273 \$6167 \$5798 \$6472 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6274 VSS \$5798 \$6167 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6275 \$6168 \$5798 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6276 \$5798 \$5798 \$6168 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6277 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6278 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6279 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6280 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6281 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6282 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6283 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6284 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6285 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6286 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6287 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6288 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6289 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6290 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6291 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6292 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6293 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6294 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6295 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6296 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6297 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6298 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6299 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6300 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6301 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6302 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6303 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6304 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6305 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6306 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6307 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6308 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6309 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6310 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6311 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6312 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6313 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6314 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6315 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6316 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6317 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6318 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6319 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6320 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6321 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6322 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6323 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6324 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6325 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6326 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6327 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6328 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6329 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6330 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6331 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6332 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6333 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6334 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6335 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6336 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6337 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6338 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6339 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6340 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6341 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6342 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6343 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6344 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6345 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6346 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6347 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6348 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6349 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6350 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6351 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6352 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6353 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6354 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6355 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6356 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6357 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6358 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6359 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6360 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6361 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6362 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6363 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6364 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6365 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6366 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6367 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6368 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6369 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6370 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6371 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6372 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6373 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6374 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6375 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6376 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6377 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6378 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6379 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6380 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6381 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6382 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6383 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6384 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6385 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6386 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6387 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6388 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6389 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6390 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6391 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6392 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6393 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6394 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6395 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6396 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6397 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6398 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6399 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6400 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6401 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6402 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6403 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6404 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6405 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6406 I1U I1U VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6407 \$7162 I1U \$7131 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6408 \$7116 I1U VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6409 \$7116 I1U \$7131 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6410 \$7162 I1U \$8504 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6411 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6412 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6413 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6414 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6415 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6416 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6417 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6418 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6419 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6420 VSS \$7132 \$7118 VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$6421 \$7118 \$7132 VSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$6422 VSS \$7132 \$7132 VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$6423 \$7132 \$7132 VSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$6424 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$6425 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$6426 VSS \$7132 \$7132 VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$6427 \$7132 \$7132 VSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$6428 VSS \$7132 \$7118 VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$6429 \$7118 \$7132 VSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$6430 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$6431 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$6432 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6433 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6434 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6435 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6436 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6437 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6438 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6439 \$7164 \$7693 \$7163 VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P
+ PS=3.62U PD=2U
M$6440 VSS \$7693 \$7164 VSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U
+ PD=3.62U
M$6441 \$7973 \$7693 \$7163 VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P
+ PS=3.62U PD=2U
M$6442 \$7974 \$7693 \$7973 VSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U
+ PD=3.62U
M$6443 \$9040 \$7693 \$7693 VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P
+ PS=3.62U PD=2U
M$6444 \$7974 \$7693 \$9040 VSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U
+ PD=3.62U
M$6445 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P PS=3.62U PD=2U
M$6446 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U PD=3.62U
M$6447 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6448 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6449 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6450 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6451 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6452 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6453 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6454 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6455 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6456 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6457 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6458 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6459 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6460 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6461 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6462 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6463 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6464 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6465 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6466 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6467 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6468 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6469 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6470 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6471 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6472 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6473 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6474 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6475 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6476 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6477 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6478 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6479 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6480 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6481 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6482 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6483 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6484 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6485 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6486 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6487 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6488 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6489 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6490 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6491 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6492 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6493 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6494 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6495 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6496 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6497 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6498 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6499 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6500 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6501 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6502 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6503 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6504 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6505 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6506 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6507 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6508 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6509 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6510 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6511 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6512 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6513 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6514 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6515 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6516 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6517 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6518 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6519 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6520 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6521 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6522 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6523 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6524 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6525 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6526 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6527 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6528 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6529 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6530 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6531 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6532 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6533 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6534 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6535 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6536 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6537 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6538 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6539 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6540 \$10111 I1U \$8504 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6541 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6542 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6543 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$6544 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$6545 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$6546 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$6547 VSS VSS VSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6548 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6549 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P PS=3.62U PD=2U
M$6550 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U PD=3.62U
M$6551 VSS VSS VSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6552 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6553 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6554 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6555 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6556 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6557 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6558 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6559 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6560 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6561 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6562 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6563 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6564 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6565 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6566 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6567 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6568 VSS \$7132 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6569 \$7081 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6570 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6571 \$7113 \$7132 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6572 VSS \$7132 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6573 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6574 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6575 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6576 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6577 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6578 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6579 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6580 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6581 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6582 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6583 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6584 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6585 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6586 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6587 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6588 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6589 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6590 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6591 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6592 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6593 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6594 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6595 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6596 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6597 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6598 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6599 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6600 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6601 \$17566 \$7693 \$7113 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6602 \$7113 \$7693 \$17566 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6603 \$17566 \$7693 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6604 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6605 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6606 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6607 \$7081 \$7693 OUT VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6608 OUT \$7693 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6609 \$7081 \$7693 OUT VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6610 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6611 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6612 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6613 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6614 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6615 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6616 \$17566 \$7693 \$7113 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6617 \$7113 \$7693 \$17566 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6618 \$17566 \$7693 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6619 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6620 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6621 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6622 OUT \$7693 \$7081 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6623 \$7081 \$7693 OUT VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6624 OUT \$7693 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6625 \$17566 \$7693 \$7113 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6626 \$7113 \$7693 \$17566 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6627 \$17566 \$7693 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6628 \$7081 \$7693 OUT VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6629 OUT \$7693 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6630 \$7081 \$7693 OUT VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6631 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6632 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6633 OUT \$7693 \$7081 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6634 \$7081 \$7693 OUT VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6635 OUT \$7693 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6636 \$17566 \$7693 \$7113 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6637 \$7113 \$7693 \$17566 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6638 \$17566 \$7693 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6639 \$7081 \$7693 OUT VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6640 OUT \$7693 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6641 \$7081 \$7693 OUT VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6642 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6643 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6644 \$17566 \$7693 \$7113 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6645 \$7113 \$7693 \$17566 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6646 \$17566 \$7693 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6647 OUT \$7693 \$7081 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6648 \$7081 \$7693 OUT VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6649 OUT \$7693 \$7081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6650 \$7113 \$7693 \$17566 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6651 \$17566 \$7693 \$7113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6652 \$7113 \$7693 \$17566 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6653 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6654 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6655 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6656 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6657 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6658 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6659 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6660 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6661 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6662 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6663 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6664 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
C$6665 \$34238 OUT 1.9208e-13 cap_mim_2f0_m4m5_noshield A=96.04P P=39.2U
C$6666 \$6 VCM 1.9208e-13 cap_mim_2f0_m4m5_noshield A=96.04P P=39.2U
C$6667 \$34238 OUT 1.9208e-13 cap_mim_2f0_m4m5_noshield A=96.04P P=39.2U
C$6668 \$6 VCM 1.9208e-13 cap_mim_2f0_m4m5_noshield A=96.04P P=39.2U
C$6669 IN_POS \$6 2e-11 cap_mim_2f0_m4m5_noshield A=10000P P=400U
C$6670 IN_POS \$6 2e-11 cap_mim_2f0_m4m5_noshield A=10000P P=400U
C$6671 IN_NEG \$34238 2e-11 cap_mim_2f0_m4m5_noshield A=10000P P=400U
C$6672 IN_NEG \$34238 2e-11 cap_mim_2f0_m4m5_noshield A=10000P P=400U
.ENDS Filter_TOP
