* Extracted by KLayout with GF180MCU LVS runset on : 16/04/2024 20:14

.SUBCKT clock_generator VSSD CK1 clks Valid VDDD OUT A B C
M$1 \$9 \$3 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$2 \$31 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$3 \$32 CK1 \$31 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$4 \$3 Valid \$32 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$5 OUT \$9 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$6 \$4 \$3 VSSD VSSD nfet_03v3 L=35U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$7 \$3 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$8 VSSD CK1 \$3 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$9 VSSD Valid \$3 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$10 \$4 \$3 \$9 VSSD nfet_03v3 L=35U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$11 \$19 \$3 VSSD VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$12 \$20 \$3 VSSD VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$13 \$21 \$3 VSSD VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$14 OUT \$9 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$15 \$19 \$3 \$33 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$16 \$20 \$3 \$34 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$17 \$21 \$3 \$35 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$18 \$9 A \$33 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$19 \$9 B \$34 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$20 \$9 C \$35 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
.ENDS clock_generator
