* Extracted by KLayout with GF180MCU LVS runset on : 29/12/2023 23:22

.SUBCKT Filter_TOP VDD A2 B2 CMOUTP CMOUTN ISBCS A1 B1 AVSS ISBCS2 IREF AVDD
+ VOUT VP VN VSS
M$1 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$4 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$5 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$6 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$7 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$8 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$9 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$10 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$11 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$12 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$13 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$14 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$15 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$16 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$17 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$18 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$19 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$20 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$21 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$22 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$23 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$24 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$25 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$26 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$27 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$28 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$29 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$30 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$31 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$32 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$33 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$34 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$35 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$36 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$37 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$38 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$39 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$40 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$41 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$42 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$43 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$44 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$45 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$46 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$47 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$48 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$49 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$50 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$51 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$52 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$53 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$54 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$55 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$56 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$57 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$58 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$59 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$60 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$61 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$62 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$63 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$64 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$65 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$66 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$67 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$68 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$69 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$70 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$71 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$72 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$73 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$74 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$75 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$76 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$77 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$78 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$79 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$80 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$81 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$82 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$83 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$84 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$85 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$86 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$87 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$88 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$89 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$90 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$91 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$92 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$93 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$94 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$95 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$96 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$97 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$98 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$99 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$100 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$101 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$102 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$103 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$104 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$105 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$106 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$107 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$108 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$109 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$110 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$111 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$112 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$113 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$114 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$115 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$116 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$117 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$118 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$119 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$120 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$121 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$122 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$123 \$136 \$173 \$917 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$124 VDD \$173 \$136 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$125 \$137 \$173 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$126 \$173 \$173 \$137 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$127 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$128 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$129 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$130 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$131 \$138 \$25 \$1 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$132 \$139 \$25 \$138 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$133 \$140 \$25 \$116 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$134 A2 \$25 \$140 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$135 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$136 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$137 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$138 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$139 \$142 \$174 \$25 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$140 \$30 \$174 \$142 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$141 \$143 \$259 \$30 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$142 \$258 \$259 \$143 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$143 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$144 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$145 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$146 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$147 \$144 \$175 \$919 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$148 VDD \$175 \$144 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$149 \$145 \$175 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$150 \$175 \$175 \$145 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$151 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$152 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$153 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$154 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$155 \$146 \$26 \$2 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$156 \$147 \$26 \$146 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$157 \$148 \$26 \$117 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$158 \$1 \$26 \$148 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$159 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$160 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$161 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$162 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$163 \$149 \$176 \$26 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$164 \$31 \$176 \$149 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$165 \$150 \$261 \$31 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$166 \$260 \$261 \$150 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$167 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$168 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$169 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$170 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$171 \$151 \$177 \$921 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$172 VDD \$177 \$151 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$173 \$152 \$177 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$174 \$177 \$177 \$152 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$175 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$176 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$177 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$178 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$179 \$153 \$27 \$3 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$180 \$154 \$27 \$153 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$181 \$155 \$27 \$118 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$182 \$2 \$27 \$155 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$183 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$184 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$185 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$186 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$187 \$156 \$178 \$27 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$188 \$32 \$178 \$156 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$189 \$157 \$263 \$32 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$190 \$262 \$263 \$157 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$191 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$192 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$193 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$194 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$195 \$158 \$179 \$923 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$196 VDD \$179 \$158 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$197 \$159 \$179 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$198 \$179 \$179 \$159 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$199 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$200 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$201 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$202 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$203 \$160 \$28 \$4 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$204 \$161 \$28 \$160 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$205 \$162 \$28 \$119 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$206 \$3 \$28 \$162 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$207 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$208 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$209 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$210 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$211 \$163 \$180 \$28 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$212 \$33 \$180 \$163 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$213 \$164 \$265 \$33 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$214 \$264 \$265 \$164 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$215 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$216 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$217 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$218 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$219 \$165 \$181 \$925 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$220 VDD \$181 \$165 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$221 \$166 \$181 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$222 \$181 \$181 \$166 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$223 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$224 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$225 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$226 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$227 \$168 \$29 B2 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$228 \$169 \$29 \$168 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$229 \$170 \$29 \$120 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$230 \$4 \$29 \$170 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$231 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$232 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$233 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$234 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$235 \$171 \$182 \$29 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$236 \$34 \$182 \$171 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$237 \$172 \$267 \$34 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$238 \$266 \$267 \$172 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$239 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$240 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$241 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$242 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$243 \$308 \$173 \$173 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$244 VDD \$173 \$308 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$245 \$309 \$173 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$246 \$917 \$173 \$309 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$247 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$248 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$249 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$250 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$251 \$310 \$25 \$174 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$252 VSS \$25 \$310 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$253 \$311 \$25 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$254 \$174 \$25 \$311 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$255 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$256 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$257 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$258 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$259 \$312 \$259 \$258 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$260 \$30 \$259 \$312 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$261 \$313 \$174 \$30 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$262 \$25 \$174 \$313 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$263 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$264 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$265 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$266 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$267 \$314 \$175 \$175 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$268 VDD \$175 \$314 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$269 \$315 \$175 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$270 \$919 \$175 \$315 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$271 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$272 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$273 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$274 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$275 \$316 \$26 \$176 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$276 VSS \$26 \$316 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$277 \$317 \$26 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$278 \$176 \$26 \$317 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$279 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$280 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$281 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$282 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$283 \$318 \$261 \$260 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$284 \$31 \$261 \$318 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$285 \$319 \$176 \$31 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$286 \$26 \$176 \$319 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$287 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$288 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$289 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$290 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$291 \$320 \$177 \$177 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$292 VDD \$177 \$320 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$293 \$321 \$177 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$294 \$921 \$177 \$321 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$295 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$296 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$297 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$298 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$299 \$322 \$27 \$178 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$300 VSS \$27 \$322 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$301 \$323 \$27 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$302 \$178 \$27 \$323 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$303 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$304 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$305 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$306 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$307 \$324 \$263 \$262 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$308 \$32 \$263 \$324 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$309 \$325 \$178 \$32 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$310 \$27 \$178 \$325 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$311 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$312 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$313 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$314 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$315 \$326 \$179 \$179 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$316 VDD \$179 \$326 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$317 \$327 \$179 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$318 \$923 \$179 \$327 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$319 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$320 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$321 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$322 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$323 \$328 \$28 \$180 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$324 VSS \$28 \$328 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$325 \$329 \$28 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$326 \$180 \$28 \$329 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$327 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$328 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$329 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$330 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$331 \$330 \$265 \$264 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$332 \$33 \$265 \$330 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$333 \$331 \$180 \$33 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$334 \$28 \$180 \$331 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$335 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$336 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$337 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$338 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$339 \$332 \$181 \$181 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$340 VDD \$181 \$332 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$341 \$333 \$181 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$342 \$925 \$181 \$333 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$343 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$344 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$345 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$346 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$347 \$334 \$29 \$182 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$348 VSS \$29 \$334 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$349 \$335 \$29 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$350 \$182 \$29 \$335 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$351 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$352 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$353 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$354 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$355 \$336 \$267 \$266 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$356 \$34 \$267 \$336 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$357 \$337 \$182 \$34 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$358 \$29 \$182 \$337 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$359 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$360 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$361 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$362 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$363 \$443 \$173 \$917 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$364 VDD \$173 \$443 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$365 \$444 \$173 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$366 \$173 \$173 \$444 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$367 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$368 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$369 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$370 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$371 \$445 \$25 \$174 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$372 VSS \$25 \$445 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$373 \$446 \$25 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$374 \$174 \$25 \$446 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$375 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$376 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$377 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$378 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$379 \$447 \$174 \$25 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$380 \$30 \$174 \$447 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$381 \$448 \$259 \$30 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$382 \$258 \$259 \$448 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$383 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$384 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$385 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$386 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$387 \$449 \$175 \$919 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$388 VDD \$175 \$449 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$389 \$450 \$175 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$390 \$175 \$175 \$450 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$391 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$392 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$393 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$394 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$395 \$451 \$26 \$176 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$396 VSS \$26 \$451 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$397 \$452 \$26 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$398 \$176 \$26 \$452 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$399 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$400 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$401 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$402 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$403 \$453 \$176 \$26 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$404 \$31 \$176 \$453 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$405 \$454 \$261 \$31 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$406 \$260 \$261 \$454 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$407 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$408 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$409 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$410 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$411 \$455 \$177 \$921 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$412 VDD \$177 \$455 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$413 \$456 \$177 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$414 \$177 \$177 \$456 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$415 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$416 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$417 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$418 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$419 \$457 \$27 \$178 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$420 VSS \$27 \$457 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$421 \$458 \$27 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$422 \$178 \$27 \$458 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$423 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$424 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$425 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$426 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$427 \$459 \$178 \$27 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$428 \$32 \$178 \$459 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$429 \$460 \$263 \$32 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$430 \$262 \$263 \$460 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$431 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$432 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$433 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$434 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$435 \$461 \$179 \$923 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$436 VDD \$179 \$461 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$437 \$462 \$179 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$438 \$179 \$179 \$462 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$439 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$440 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$441 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$442 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$443 \$463 \$28 \$180 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$444 VSS \$28 \$463 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$445 \$464 \$28 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$446 \$180 \$28 \$464 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$447 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$448 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$449 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$450 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$451 \$465 \$180 \$28 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$452 \$33 \$180 \$465 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$453 \$466 \$265 \$33 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$454 \$264 \$265 \$466 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$455 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$456 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$457 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$458 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$459 \$467 \$181 \$925 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$460 VDD \$181 \$467 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$461 \$468 \$181 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$462 \$181 \$181 \$468 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$463 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$464 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$465 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$466 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$467 \$469 \$29 \$182 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$468 VSS \$29 \$469 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$469 \$470 \$29 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$470 \$182 \$29 \$470 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$471 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$472 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$473 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$474 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$475 \$471 \$182 \$29 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$476 \$34 \$182 \$471 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$477 \$472 \$267 \$34 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$478 \$266 \$267 \$472 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$479 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$480 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$481 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$482 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$483 \$588 \$173 \$173 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$484 VDD \$173 \$588 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$485 \$589 \$173 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$486 \$917 \$173 \$589 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$487 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$488 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$489 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$490 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$491 \$590 \$25 A2 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$492 \$116 \$25 \$590 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$493 \$591 \$25 \$139 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$494 \$1 \$25 \$591 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$495 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$496 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$497 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$498 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$499 \$592 \$259 \$258 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$500 \$30 \$259 \$592 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$501 \$593 \$174 \$30 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$502 \$25 \$174 \$593 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$503 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$504 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$505 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$506 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$507 \$594 \$175 \$175 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$508 VDD \$175 \$594 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$509 \$595 \$175 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$510 \$919 \$175 \$595 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$511 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$512 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$513 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$514 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$515 \$596 \$26 \$1 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$516 \$117 \$26 \$596 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$517 \$597 \$26 \$147 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$518 \$2 \$26 \$597 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$519 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$520 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$521 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$522 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$523 \$598 \$261 \$260 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$524 \$31 \$261 \$598 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$525 \$599 \$176 \$31 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$526 \$26 \$176 \$599 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$527 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$528 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$529 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$530 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$531 \$600 \$177 \$177 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$532 VDD \$177 \$600 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$533 \$601 \$177 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$534 \$921 \$177 \$601 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$535 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$536 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$537 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$538 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$539 \$602 \$27 \$2 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$540 \$118 \$27 \$602 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$541 \$603 \$27 \$154 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$542 \$3 \$27 \$603 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$543 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$544 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$545 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$546 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$547 \$604 \$263 \$262 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$548 \$32 \$263 \$604 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$549 \$605 \$178 \$32 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$550 \$27 \$178 \$605 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$551 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$552 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$553 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$554 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$555 \$606 \$179 \$179 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$556 VDD \$179 \$606 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$557 \$607 \$179 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$558 \$923 \$179 \$607 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$559 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$560 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$561 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$562 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$563 \$608 \$28 \$3 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$564 \$119 \$28 \$608 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$565 \$609 \$28 \$161 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$566 \$4 \$28 \$609 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$567 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$568 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$569 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$570 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$571 \$610 \$265 \$264 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$572 \$33 \$265 \$610 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$573 \$611 \$180 \$33 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$574 \$28 \$180 \$611 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$575 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$576 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$577 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$578 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$579 \$612 \$181 \$181 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$580 VDD \$181 \$612 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$581 \$613 \$181 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$582 \$925 \$181 \$613 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$583 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$584 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$585 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$586 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$587 \$614 \$29 \$4 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$588 \$120 \$29 \$614 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$589 \$615 \$29 \$169 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$590 B2 \$29 \$615 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$591 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$592 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$593 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$594 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$595 \$616 \$267 \$266 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$596 \$34 \$267 \$616 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$597 \$617 \$182 \$34 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$598 \$29 \$182 \$617 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$599 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$600 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$601 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$602 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$603 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$604 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$605 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$606 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$607 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$608 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$609 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$610 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$611 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$612 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$613 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$614 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$615 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$616 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$617 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$618 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$619 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$620 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$621 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$622 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$623 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$624 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$625 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$626 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$627 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$628 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$629 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$630 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$631 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$632 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$633 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$634 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$635 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$636 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$637 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$638 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$639 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$640 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$641 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$642 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$643 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$644 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$645 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$646 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$647 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$648 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$649 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$650 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$651 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$652 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$653 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$654 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$655 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$656 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$657 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$658 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$659 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$660 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$661 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$662 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$663 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$664 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$665 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$666 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$667 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$668 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$669 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$670 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$671 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$672 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$673 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$674 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$675 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$676 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$677 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$678 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$679 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$680 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$681 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$682 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$683 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$684 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$685 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$686 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$687 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$688 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$689 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$690 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$691 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$692 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$693 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$694 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$695 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$696 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$697 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$698 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$699 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$700 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$701 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$702 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$703 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$704 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$705 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$706 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$707 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$708 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$709 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$710 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$711 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$712 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$713 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$714 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$715 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$716 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$717 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$718 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$719 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$720 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$721 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$722 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$723 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$724 \$1583 \$1573 \$1582 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$725 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$726 \$1670 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$727 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$728 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$729 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$730 \$1584 \$1573 \$1583 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$731 \$1585 \$1573 \$1584 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$732 \$1586 \$1573 \$1585 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$733 \$1671 \$1573 \$1670 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$734 \$1672 \$1573 \$1671 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$735 \$1673 \$1573 \$1672 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$736 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$737 VDD \$1573 \$1586 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$738 \$1674 \$1573 \$1673 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$739 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$740 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$741 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$742 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$743 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$744 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$745 \$1675 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$746 \$1588 \$1573 \$1587 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$747 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$748 \$1589 \$1573 \$1588 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$749 \$1590 \$1573 \$1589 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$750 \$1591 \$1573 \$1590 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$751 \$1676 \$1573 \$1675 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$752 \$1677 \$1573 \$1676 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$753 \$1678 \$1573 \$1677 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$754 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$755 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$756 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$757 VDD \$1573 \$1591 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$758 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$759 \$1679 \$1573 \$1678 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$760 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$761 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$762 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$763 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$764 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$765 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$766 \$1680 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$767 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$768 \$1593 \$1573 \$1592 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$769 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$770 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$771 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$772 \$1594 \$1573 \$1593 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$773 \$1595 \$1573 \$1594 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$774 \$1596 \$1573 \$1595 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$775 \$1681 \$1573 \$1680 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$776 \$1682 \$1573 \$1681 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$777 \$1683 \$1573 \$1682 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$778 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$779 VDD \$1573 \$1596 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$780 \$1684 \$1573 \$1683 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$781 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$782 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$783 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$784 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$785 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$786 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$787 \$1685 \$1574 \$174 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$788 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$789 \$1598 \$1574 \$1597 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$790 \$1686 \$1574 \$1685 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$791 \$1687 \$1574 \$1686 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$792 \$1688 \$1574 \$1687 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$793 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$794 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$795 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$796 \$1599 \$1574 \$1598 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$797 \$1600 \$1574 \$1599 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$798 \$1601 \$1574 \$1600 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$799 \$1602 \$1574 \$1601 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$800 \$1689 \$1574 \$1688 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$801 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$802 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$803 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$804 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$805 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$806 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$807 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$808 \$1690 \$1574 \$176 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$809 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$810 \$1604 \$1574 \$1603 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$811 \$1605 \$1574 \$1604 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$812 \$1606 \$1574 \$1605 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$813 \$1607 \$1574 \$1606 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$814 \$1691 \$1574 \$1690 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$815 \$1692 \$1574 \$1691 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$816 \$1693 \$1574 \$1692 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$817 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$818 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$819 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$820 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$821 \$1608 \$1574 \$1607 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$822 \$1694 \$1574 \$1693 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$823 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$824 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$825 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$826 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$827 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$828 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$829 \$1610 \$1574 \$1609 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$830 \$1695 \$1574 \$178 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$831 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$832 \$1696 \$1574 \$1695 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$833 \$1697 \$1574 \$1696 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$834 \$1698 \$1574 \$1697 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$835 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$836 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$837 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$838 \$1611 \$1574 \$1610 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$839 \$1612 \$1574 \$1611 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$840 \$1613 \$1574 \$1612 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$841 \$1699 \$1574 \$1698 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$842 \$1614 \$1574 \$1613 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$843 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$844 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$845 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$846 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$847 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$848 \$1820 \$1573 \$1819 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$849 \$1821 \$1573 \$1820 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$850 \$1822 \$1573 \$1821 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$851 \$1823 \$1573 \$1822 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$852 \$1674 \$1573 \$1823 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$853 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$854 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$855 \$1825 \$1573 \$1824 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$856 \$1826 \$1573 \$1825 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$857 \$1827 \$1573 \$1826 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$858 \$1828 \$1573 \$1827 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$859 \$1679 \$1573 \$1828 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$860 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$861 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$862 \$1830 \$1573 \$1829 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$863 \$1831 \$1573 \$1830 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$864 \$1832 \$1573 \$1831 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$865 \$1833 \$1573 \$1832 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$866 \$1684 \$1573 \$1833 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$867 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$868 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$869 \$1835 \$1574 \$1834 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$870 \$1836 \$1574 \$1835 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$871 \$1837 \$1574 \$1836 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$872 \$1838 \$1574 \$1837 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$873 \$1689 \$1574 \$1838 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$874 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$875 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$876 \$1840 \$1574 \$1839 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$877 \$1841 \$1574 \$1840 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$878 \$1842 \$1574 \$1841 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$879 \$1843 \$1574 \$1842 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$880 \$1694 \$1574 \$1843 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$881 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$882 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$883 \$1845 \$1574 \$1844 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$884 \$1846 \$1574 \$1845 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$885 \$1847 \$1574 \$1846 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$886 \$1848 \$1574 \$1847 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$887 \$1699 \$1574 \$1848 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$888 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$889 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$890 \$1975 \$1573 \$1819 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$891 \$1976 \$1573 \$1975 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$892 \$1977 \$1573 \$1976 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$893 \$1978 \$1573 \$1977 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$894 \$1979 \$1573 \$1978 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$895 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$896 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$897 \$1980 \$1573 \$1824 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$898 \$1981 \$1573 \$1980 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$899 \$1982 \$1573 \$1981 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$900 \$1983 \$1573 \$1982 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$901 \$1984 \$1573 \$1983 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$902 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$903 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$904 \$1985 \$1573 \$1829 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$905 \$1986 \$1573 \$1985 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$906 \$1987 \$1573 \$1986 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$907 \$1988 \$1573 \$1987 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$908 \$1989 \$1573 \$1988 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$909 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$910 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$911 \$1990 \$1574 \$1834 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$912 \$1991 \$1574 \$1990 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$913 \$1992 \$1574 \$1991 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$914 \$1993 \$1574 \$1992 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$915 \$1994 \$1574 \$1993 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$916 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$917 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$918 \$1995 \$1574 \$1839 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$919 \$1996 \$1574 \$1995 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$920 \$1997 \$1574 \$1996 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$921 \$1998 \$1574 \$1997 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$922 \$1999 \$1574 \$1998 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$923 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$924 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$925 \$2000 \$1574 \$1844 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$926 \$2001 \$1574 \$2000 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$927 \$2002 \$1574 \$2001 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$928 \$2003 \$1574 \$2002 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$929 \$2004 \$1574 \$2003 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$930 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$931 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$932 \$2146 \$1573 \$1582 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$933 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$934 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$935 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$936 \$2148 \$1573 \$2147 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$937 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$938 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$939 \$2149 \$1573 \$1587 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$940 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$941 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$942 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$943 \$2151 \$1573 \$2150 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$944 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$945 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$946 \$2152 \$1573 \$1592 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$947 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$948 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$949 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$950 \$2153 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$951 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$952 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$953 \$2154 \$1574 \$1597 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$954 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$955 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$956 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$957 \$2155 \$1574 \$1602 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$958 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$959 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$960 \$2156 \$1574 \$1603 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$961 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$962 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$963 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$964 \$2157 \$1574 \$1608 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$965 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$966 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$967 \$2158 \$1574 \$1609 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$968 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$969 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$970 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$971 \$2159 \$1574 \$1614 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$972 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$973 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$974 \$2146 \$1573 \$2289 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$975 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$976 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$977 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$978 \$2148 \$1573 \$2290 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$979 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$980 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$981 \$2149 \$1573 \$2291 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$982 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$983 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$984 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$985 \$2151 \$1573 \$2292 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$986 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$987 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$988 \$2152 \$1573 \$2293 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$989 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$990 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$991 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$992 \$2153 \$1573 \$2294 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$993 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$994 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$995 \$2154 \$1574 \$2295 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$996 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$997 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$998 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$999 \$2155 \$1574 \$30 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1000 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1001 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1002 \$2156 \$1574 \$2296 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1003 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1004 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1005 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1006 \$2157 \$1574 \$31 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1007 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1008 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1009 \$2158 \$1574 \$2297 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1010 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1011 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1012 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1013 \$2159 \$1574 \$32 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1014 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1015 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1016 \$2446 \$1573 \$2445 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1017 \$2447 \$1573 \$2446 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1018 \$2448 \$1573 \$2447 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1019 \$2449 \$1573 \$2448 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1020 \$1979 \$1573 \$2449 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1021 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1022 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1023 \$2451 \$1573 \$2450 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1024 \$2452 \$1573 \$2451 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1025 \$2453 \$1573 \$2452 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1026 \$2454 \$1573 \$2453 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1027 \$1984 \$1573 \$2454 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1028 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1029 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1030 \$2456 \$1573 \$2455 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1031 \$2457 \$1573 \$2456 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1032 \$2458 \$1573 \$2457 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1033 \$2459 \$1573 \$2458 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1034 \$1989 \$1573 \$2459 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1035 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1036 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1037 \$2461 \$1574 \$2460 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1038 \$2462 \$1574 \$2461 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1039 \$2463 \$1574 \$2462 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1040 \$2464 \$1574 \$2463 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1041 \$1994 \$1574 \$2464 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1042 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1043 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1044 \$2466 \$1574 \$2465 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1045 \$2467 \$1574 \$2466 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1046 \$2468 \$1574 \$2467 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1047 \$2469 \$1574 \$2468 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1048 \$1999 \$1574 \$2469 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1049 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1050 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1051 \$2471 \$1574 \$2470 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1052 \$2472 \$1574 \$2471 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1053 \$2473 \$1574 \$2472 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1054 \$2474 \$1574 \$2473 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1055 \$2004 \$1574 \$2474 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1056 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1057 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1058 \$2619 \$1573 \$2445 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1059 \$2620 \$1573 \$2619 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1060 \$2621 \$1573 \$2620 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1061 \$2622 \$1573 \$2621 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1062 \$2623 \$1573 \$2622 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1063 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1064 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1065 \$2624 \$1573 \$2450 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1066 \$2625 \$1573 \$2624 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1067 \$2626 \$1573 \$2625 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1068 \$2627 \$1573 \$2626 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1069 \$2628 \$1573 \$2627 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1070 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1071 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1072 \$2629 \$1573 \$2455 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1073 \$2630 \$1573 \$2629 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1074 \$2631 \$1573 \$2630 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1075 \$2632 \$1573 \$2631 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1076 \$2633 \$1573 \$2632 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1077 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1078 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1079 \$2634 \$1574 \$2460 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1080 \$2635 \$1574 \$2634 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1081 \$2636 \$1574 \$2635 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1082 \$2637 \$1574 \$2636 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1083 \$2638 \$1574 \$2637 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1084 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1085 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1086 \$2639 \$1574 \$2465 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1087 \$2640 \$1574 \$2639 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1088 \$2641 \$1574 \$2640 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1089 \$2642 \$1574 \$2641 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1090 \$2643 \$1574 \$2642 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1091 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1092 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1093 \$2644 \$1574 \$2470 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1094 \$2645 \$1574 \$2644 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1095 \$2646 \$1574 \$2645 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1096 \$2647 \$1574 \$2646 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1097 \$2648 \$1574 \$2647 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1098 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1099 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1100 \$2787 \$1573 \$5958 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1101 \$2788 \$1573 \$2787 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1102 \$2789 \$1573 \$2788 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1103 \$2790 \$1573 \$2789 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1104 \$2623 \$1573 \$2790 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1105 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1106 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1107 \$2791 \$1573 \$5959 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1108 \$2792 \$1573 \$2791 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1109 \$2793 \$1573 \$2792 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1110 \$2794 \$1573 \$2793 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1111 \$2628 \$1573 \$2794 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1112 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1113 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1114 \$2796 \$1573 CMOUTP VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1115 \$2797 \$1573 \$2796 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1116 \$2798 \$1573 \$2797 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1117 \$2799 \$1573 \$2798 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1118 \$2633 \$1573 \$2799 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1119 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1120 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1121 \$2800 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1122 \$2801 \$1574 \$2800 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1123 \$2802 \$1574 \$2801 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1124 \$2803 \$1574 \$2802 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1125 \$2638 \$1574 \$2803 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1126 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1127 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1128 \$2804 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1129 \$2805 \$1574 \$2804 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1130 \$2806 \$1574 \$2805 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1131 \$2807 \$1574 \$2806 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1132 \$2643 \$1574 \$2807 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1133 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1134 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1135 \$2808 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1136 \$2809 \$1574 \$2808 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1137 \$2810 \$1574 \$2809 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1138 \$2811 \$1574 \$2810 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1139 \$2648 \$1574 \$2811 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1140 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1141 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1142 \$2941 \$1573 \$2289 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1143 \$2942 \$1573 \$2941 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1144 \$2943 \$1573 \$2942 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1145 \$2944 \$1573 \$2943 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1146 \$2290 \$1573 \$2944 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1147 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1148 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1149 \$2945 \$1573 \$2291 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1150 \$2946 \$1573 \$2945 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1151 \$2947 \$1573 \$2946 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1152 \$2948 \$1573 \$2947 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1153 \$2292 \$1573 \$2948 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1154 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1155 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1156 \$2949 \$1573 \$2293 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1157 \$2950 \$1573 \$2949 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1158 \$2951 \$1573 \$2950 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1159 \$2952 \$1573 \$2951 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1160 \$2294 \$1573 \$2952 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1161 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1162 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1163 \$2953 \$1574 \$2295 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1164 \$2954 \$1574 \$2953 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1165 \$2955 \$1574 \$2954 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1166 \$2956 \$1574 \$2955 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1167 VDD \$1574 \$2956 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1168 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1169 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1170 \$2957 \$1574 \$2296 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1171 \$2958 \$1574 \$2957 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1172 \$2959 \$1574 \$2958 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1173 \$2960 \$1574 \$2959 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1174 VDD \$1574 \$2960 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1175 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1176 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1177 \$2961 \$1574 \$2297 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1178 \$2962 \$1574 \$2961 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1179 \$2963 \$1574 \$2962 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1180 \$2964 \$1574 \$2963 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1181 VDD \$1574 \$2964 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1182 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1183 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1184 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1185 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1186 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1187 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1188 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1189 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1190 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1191 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1192 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1193 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1194 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1195 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1196 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1197 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1198 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1199 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1200 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1201 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1202 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1203 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1204 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1205 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1206 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1207 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1208 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1209 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1210 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1211 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1212 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1213 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1214 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1215 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1216 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1217 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1218 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1219 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1220 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1221 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1222 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1223 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1224 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1225 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1226 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1227 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1228 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1229 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1230 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1231 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1232 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1233 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1234 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1235 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1236 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1237 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1238 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1239 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1240 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1241 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1242 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1243 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1244 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1245 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1246 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1247 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1248 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1249 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1250 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1251 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1252 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1253 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1254 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1255 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1256 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1257 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1258 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1259 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1260 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1261 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1262 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1263 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1264 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1265 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1266 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1267 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1268 \$3266 \$1573 \$3265 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1269 \$3267 \$1573 \$3266 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1270 \$3268 \$1573 \$3267 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1271 \$3269 \$1573 \$3268 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1272 VDD \$1573 \$3269 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1273 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1274 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1275 \$3271 \$1573 \$3270 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1276 \$3272 \$1573 \$3271 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1277 \$3273 \$1573 \$3272 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1278 \$3274 \$1573 \$3273 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1279 VDD \$1573 \$3274 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1280 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1281 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1282 \$3276 \$1573 \$3275 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1283 \$3277 \$1573 \$3276 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1284 \$3278 \$1573 \$3277 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1285 \$3279 \$1573 \$3278 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1286 VDD \$1573 \$3279 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1287 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1288 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1289 \$3281 \$1574 \$3280 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1290 \$3282 \$1574 \$3281 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1291 \$3283 \$1574 \$3282 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1292 \$3284 \$1574 \$3283 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1293 \$3285 \$1574 \$3284 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1294 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1295 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1296 \$3287 \$1574 \$3286 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1297 \$3288 \$1574 \$3287 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1298 \$3289 \$1574 \$3288 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1299 \$3290 \$1574 \$3289 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1300 \$3291 \$1574 \$3290 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1301 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1302 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1303 \$3293 \$1574 \$3292 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1304 \$3294 \$1574 \$3293 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1305 \$3295 \$1574 \$3294 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1306 \$3296 \$1574 \$3295 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1307 \$3297 \$1574 \$3296 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1308 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1309 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1310 \$3440 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1311 \$3441 \$1573 \$3440 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1312 \$3442 \$1573 \$3441 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1313 \$3443 \$1573 \$3442 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1314 \$3444 \$1573 \$3443 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1315 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1316 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1317 \$3445 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1318 \$3446 \$1573 \$3445 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1319 \$3447 \$1573 \$3446 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1320 \$3448 \$1573 \$3447 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1321 \$3449 \$1573 \$3448 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1322 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1323 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1324 \$3450 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1325 \$3451 \$1573 \$3450 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1326 \$3452 \$1573 \$3451 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1327 \$3453 \$1573 \$3452 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1328 \$3454 \$1573 \$3453 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1329 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1330 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1331 \$3455 \$1574 \$180 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1332 \$3456 \$1574 \$3455 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1333 \$3457 \$1574 \$3456 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1334 \$3458 \$1574 \$3457 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1335 \$3459 \$1574 \$3458 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1336 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1337 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1338 \$3460 \$1574 \$182 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1339 \$3461 \$1574 \$3460 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1340 \$3462 \$1574 \$3461 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1341 \$3463 \$1574 \$3462 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1342 \$3464 \$1574 \$3463 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1343 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1344 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1345 \$3465 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1346 \$3466 \$1574 \$3465 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1347 \$3467 \$1574 \$3466 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1348 \$3468 \$1574 \$3467 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1349 \$3469 \$1574 \$3468 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1350 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1351 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1352 \$3606 \$1573 \$3605 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1353 \$3607 \$1573 \$3606 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1354 \$3608 \$1573 \$3607 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1355 \$3609 \$1573 \$3608 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1356 \$3444 \$1573 \$3609 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1357 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1358 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1359 \$3611 \$1573 \$3610 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1360 \$3612 \$1573 \$3611 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1361 \$3613 \$1573 \$3612 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1362 \$3614 \$1573 \$3613 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1363 \$3449 \$1573 \$3614 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1364 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1365 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1366 \$3616 \$1573 \$3615 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1367 \$3617 \$1573 \$3616 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1368 \$3618 \$1573 \$3617 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1369 \$3619 \$1573 \$3618 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1370 \$3454 \$1573 \$3619 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1371 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1372 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1373 \$3621 \$1574 \$3620 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1374 \$3622 \$1574 \$3621 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1375 \$3623 \$1574 \$3622 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1376 \$3624 \$1574 \$3623 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1377 \$3459 \$1574 \$3624 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1378 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1379 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1380 \$3626 \$1574 \$3625 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1381 \$3627 \$1574 \$3626 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1382 \$3628 \$1574 \$3627 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1383 \$3629 \$1574 \$3628 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1384 \$3464 \$1574 \$3629 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1385 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1386 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1387 \$3631 \$1574 \$3630 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1388 \$3632 \$1574 \$3631 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1389 \$3633 \$1574 \$3632 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1390 \$3634 \$1574 \$3633 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1391 \$3469 \$1574 \$3634 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1392 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1393 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1394 \$3761 \$1573 \$3605 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1395 \$3762 \$1573 \$3761 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1396 \$3763 \$1573 \$3762 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1397 \$3764 \$1573 \$3763 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1398 \$3765 \$1573 \$3764 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1399 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1400 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1401 \$3766 \$1573 \$3610 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1402 \$3767 \$1573 \$3766 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1403 \$3768 \$1573 \$3767 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1404 \$3769 \$1573 \$3768 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1405 \$3770 \$1573 \$3769 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1406 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1407 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1408 \$3771 \$1573 \$3615 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1409 \$3772 \$1573 \$3771 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1410 \$3773 \$1573 \$3772 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1411 \$3774 \$1573 \$3773 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1412 \$3775 \$1573 \$3774 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1413 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1414 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1415 \$3776 \$1574 \$3620 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1416 \$3777 \$1574 \$3776 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1417 \$3778 \$1574 \$3777 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1418 \$3779 \$1574 \$3778 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1419 \$3780 \$1574 \$3779 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1420 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1421 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1422 \$3781 \$1574 \$3625 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1423 \$3782 \$1574 \$3781 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1424 \$3783 \$1574 \$3782 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1425 \$3784 \$1574 \$3783 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1426 \$3785 \$1574 \$3784 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1427 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1428 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1429 \$3786 \$1574 \$3630 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1430 \$3787 \$1574 \$3786 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1431 \$3788 \$1574 \$3787 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1432 \$3789 \$1574 \$3788 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1433 \$3790 \$1574 \$3789 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1434 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1435 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1436 \$3925 \$1573 \$3265 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1437 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1438 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1439 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1440 \$3926 \$1573 \$3943 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1441 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1442 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1443 \$3927 \$1573 \$3270 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1444 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1445 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1446 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1447 \$3928 \$1573 \$3944 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1448 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1449 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1450 \$3929 \$1573 \$3275 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1451 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1452 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1453 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1454 \$3930 \$1573 \$3945 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1455 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1456 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1457 \$3931 \$1574 \$3280 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1458 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1459 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1460 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1461 \$3932 \$1574 \$3285 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1462 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1463 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1464 \$3933 \$1574 \$3286 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1465 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1466 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1467 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1468 \$3934 \$1574 \$3291 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1469 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1470 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1471 \$3935 \$1574 \$3292 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1472 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1473 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1474 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1475 \$3936 \$1574 \$3297 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1476 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1477 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1478 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1479 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1480 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1481 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1482 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1483 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1484 \$3925 \$1573 \$4094 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1485 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1486 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1487 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1488 \$3926 \$1573 \$4095 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1489 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1490 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1491 \$3927 \$1573 \$4096 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1492 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1493 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1494 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1495 \$3928 \$1573 \$4097 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1496 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1497 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1498 \$3929 \$1573 \$4098 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1499 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1500 \$1573 \$1573 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1501 VDD \$1573 \$1573 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1502 \$3930 \$1573 \$4099 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1503 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1504 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1505 \$3931 \$1574 \$4100 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1506 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1507 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1508 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1509 \$3932 \$1574 \$33 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1510 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1511 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1512 \$3933 \$1574 \$4101 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1513 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1514 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1515 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1516 \$3934 \$1574 \$34 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1517 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1518 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1519 \$3935 \$1574 \$4102 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1520 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1521 VDD \$1574 \$1574 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1522 \$1574 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1523 \$3936 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1524 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1525 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1526 \$4158 \$4093 \$1773 VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1527 VDD \$4093 \$4158 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1528 \$4159 \$4093 VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1529 \$1730 \$4093 \$4159 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1530 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1531 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1532 \$4262 \$1573 \$4261 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1533 \$4263 \$1573 \$4262 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1534 \$4264 \$1573 \$4263 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1535 \$4265 \$1573 \$4264 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1536 \$3765 \$1573 \$4265 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1537 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1538 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1539 \$4267 \$1573 \$4266 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1540 \$4268 \$1573 \$4267 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1541 \$4269 \$1573 \$4268 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1542 \$4270 \$1573 \$4269 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1543 \$3770 \$1573 \$4270 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1544 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1545 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1546 \$4272 \$1573 \$4271 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1547 \$4273 \$1573 \$4272 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1548 \$4274 \$1573 \$4273 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1549 \$4275 \$1573 \$4274 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1550 \$3775 \$1573 \$4275 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1551 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1552 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1553 \$4277 \$1574 \$4276 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1554 \$4278 \$1574 \$4277 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1555 \$4279 \$1574 \$4278 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1556 \$4280 \$1574 \$4279 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1557 \$3780 \$1574 \$4280 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1558 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1559 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1560 \$4282 \$1574 \$4281 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1561 \$4283 \$1574 \$4282 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1562 \$4284 \$1574 \$4283 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1563 \$4285 \$1574 \$4284 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1564 \$3785 \$1574 \$4285 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1565 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1566 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1567 \$4287 \$1574 \$4286 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1568 \$4288 \$1574 \$4287 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1569 \$4289 \$1574 \$4288 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1570 \$4290 \$1574 \$4289 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1571 \$3790 \$1574 \$4290 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1572 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1573 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1574 \$4341 \$4093 \$4093 VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1575 VDD \$4093 \$4341 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1576 \$4342 \$4093 VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1577 \$4093 \$4093 \$4342 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1578 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1579 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1580 \$4444 \$1573 \$4261 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1581 \$4445 \$1573 \$4444 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1582 \$4446 \$1573 \$4445 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1583 \$4447 \$1573 \$4446 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1584 \$4448 \$1573 \$4447 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1585 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1586 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1587 \$4449 \$1573 \$4266 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1588 \$4450 \$1573 \$4449 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1589 \$4451 \$1573 \$4450 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1590 \$4452 \$1573 \$4451 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1591 \$4453 \$1573 \$4452 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1592 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1593 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1594 \$4454 \$1573 \$4271 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1595 \$4455 \$1573 \$4454 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1596 \$4456 \$1573 \$4455 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1597 \$4457 \$1573 \$4456 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1598 \$4458 \$1573 \$4457 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1599 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1600 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1601 \$4459 \$1574 \$4276 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1602 \$4460 \$1574 \$4459 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1603 \$4461 \$1574 \$4460 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1604 \$4462 \$1574 \$4461 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1605 \$4463 \$1574 \$4462 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1606 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1607 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1608 \$4464 \$1574 \$4281 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1609 \$4465 \$1574 \$4464 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1610 \$4466 \$1574 \$4465 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1611 \$4467 \$1574 \$4466 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1612 \$4468 \$1574 \$4467 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1613 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1614 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1615 \$4469 \$1574 \$4286 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1616 \$4470 \$1574 \$4469 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1617 \$4471 \$1574 \$4470 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1618 \$4472 \$1574 \$4471 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1619 \$4473 \$1574 \$4472 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1620 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1621 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1622 \$4515 \$4093 \$1730 VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1623 VDD \$4093 \$4515 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1624 \$4516 \$4093 VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1625 \$1773 \$4093 \$4516 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1626 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1627 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1628 \$4608 \$1573 \$5955 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1629 \$4609 \$1573 \$4608 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1630 \$4610 \$1573 \$4609 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1631 \$4611 \$1573 \$4610 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1632 \$4448 \$1573 \$4611 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1633 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1634 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1635 \$4612 \$1573 \$5956 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1636 \$4613 \$1573 \$4612 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1637 \$4614 \$1573 \$4613 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1638 \$4615 \$1573 \$4614 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1639 \$4453 \$1573 \$4615 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1640 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1641 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1642 \$4616 \$1573 \$5957 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1643 \$4617 \$1573 \$4616 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1644 \$4618 \$1573 \$4617 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1645 \$4619 \$1573 \$4618 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1646 \$4458 \$1573 \$4619 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1647 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1648 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1649 \$4620 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1650 \$4621 \$1574 \$4620 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1651 \$4622 \$1574 \$4621 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1652 \$4623 \$1574 \$4622 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1653 \$4463 \$1574 \$4623 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1654 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1655 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1656 \$4624 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1657 \$4625 \$1574 \$4624 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1658 \$4626 \$1574 \$4625 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1659 \$4627 \$1574 \$4626 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1660 \$4468 \$1574 \$4627 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1661 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1662 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1663 \$4628 \$1574 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1664 \$4629 \$1574 \$4628 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1665 \$4630 \$1574 \$4629 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1666 \$4631 \$1574 \$4630 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1667 \$4473 \$1574 \$4631 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1668 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1669 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1670 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1671 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1672 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1673 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1674 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1675 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1676 \$4756 \$1573 \$4094 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1677 \$4757 \$1573 \$4756 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1678 \$4758 \$1573 \$4757 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1679 \$4759 \$1573 \$4758 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1680 \$4095 \$1573 \$4759 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1681 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1682 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1683 \$4760 \$1573 \$4096 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1684 \$4761 \$1573 \$4760 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1685 \$4762 \$1573 \$4761 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1686 \$4763 \$1573 \$4762 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1687 \$4097 \$1573 \$4763 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1688 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1689 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1690 \$4764 \$1573 \$4098 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1691 \$4765 \$1573 \$4764 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1692 \$4766 \$1573 \$4765 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1693 \$4767 \$1573 \$4766 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1694 \$4099 \$1573 \$4767 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1695 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1696 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1697 \$4768 \$1574 \$4100 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1698 \$4769 \$1574 \$4768 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1699 \$4770 \$1574 \$4769 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1700 \$4771 \$1574 \$4770 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1701 VDD \$1574 \$4771 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1702 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1703 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1704 \$4772 \$1574 \$4101 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1705 \$4773 \$1574 \$4772 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1706 \$4774 \$1574 \$4773 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1707 \$4775 \$1574 \$4774 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1708 VDD \$1574 \$4775 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1709 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1710 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1711 \$4776 \$1574 \$4102 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U
+ PD=5.3U
M$1712 \$4777 \$1574 \$4776 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1713 \$4778 \$1574 \$4777 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1714 \$4779 \$1574 \$4778 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1715 VDD \$1574 \$4779 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1716 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1717 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1718 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1719 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1720 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1721 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1722 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1723 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1724 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1725 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1726 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1727 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1728 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1729 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1730 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1731 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1732 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1733 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1734 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1735 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1736 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1737 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1738 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1739 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1740 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1741 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1742 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1743 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1744 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1745 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1746 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1747 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1748 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1749 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1750 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1751 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1752 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1753 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1754 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1755 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$1756 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1757 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1758 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1759 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1760 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1761 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1762 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1763 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1764 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1765 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1766 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1767 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1768 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1769 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1770 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1771 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1772 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1773 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1774 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1775 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1776 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1777 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1778 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1779 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1780 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1781 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1782 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1783 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1784 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1785 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1786 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1787 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1788 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1789 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1790 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1791 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1792 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1793 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1794 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1795 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1796 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1797 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1798 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1799 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1800 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1801 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1802 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1803 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1804 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1805 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1806 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1807 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1808 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1809 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1810 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1811 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1812 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1813 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1814 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1815 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1816 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1817 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1818 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1819 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1820 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1821 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1822 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1823 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1824 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1825 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1826 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1827 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1828 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1829 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1830 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1831 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1832 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1833 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1834 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1835 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1836 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1837 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1838 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1839 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1840 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1841 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1842 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1843 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1844 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1845 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1846 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1847 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1848 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1849 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1850 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1851 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1852 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1853 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1854 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1855 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1856 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1857 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1858 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1859 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1860 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1861 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1862 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1863 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1864 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1865 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1866 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1867 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1868 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1869 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1870 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1871 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1872 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1873 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1874 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1875 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1876 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1877 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1878 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1879 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1880 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1881 \$5814 \$5073 \$5073 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1882 VDD \$5073 \$5814 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1883 \$5815 \$5073 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1884 \$4973 \$5073 \$5815 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1885 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1886 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1887 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1888 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1889 \$5817 \$5850 A1 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1890 \$5076 \$5850 \$5817 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1891 \$5818 \$5850 \$5183 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1892 \$5819 \$5850 \$5818 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1893 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1894 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1895 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1896 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1897 \$5820 \$5113 \$5114 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1898 \$3943 \$5113 \$5820 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1899 \$5821 \$5955 \$3943 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1900 \$5850 \$5955 \$5821 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1901 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1902 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1903 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1904 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1905 \$5822 \$5081 \$5081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1906 VDD \$5081 \$5822 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1907 \$5823 \$5081 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1908 \$4974 \$5081 \$5823 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1909 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1910 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1911 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1912 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1913 \$5824 \$5851 \$5819 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1914 \$5084 \$5851 \$5824 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1915 \$5825 \$5851 \$5184 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1916 \$5826 \$5851 \$5825 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1917 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1918 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1919 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1920 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1921 \$5827 \$5115 \$5116 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1922 \$3944 \$5115 \$5827 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1923 \$5828 \$5956 \$3944 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1924 \$5851 \$5956 \$5828 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1925 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1926 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1927 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1928 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1929 \$5829 \$5089 \$5089 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1930 VDD \$5089 \$5829 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1931 \$5830 \$5089 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1932 \$4975 \$5089 \$5830 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1933 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1934 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1935 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1936 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1937 \$5831 \$5852 \$5826 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1938 \$5092 \$5852 \$5831 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1939 \$5832 \$5852 \$5185 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1940 \$5833 \$5852 \$5832 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1941 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1942 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1943 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1944 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1945 \$5834 \$5117 \$5118 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1946 \$3945 \$5117 \$5834 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1947 \$5835 \$5957 \$3945 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1948 \$5852 \$5957 \$5835 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1949 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1950 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1951 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1952 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1953 \$5836 \$5097 \$5097 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1954 VDD \$5097 \$5836 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1955 \$5837 \$5097 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1956 \$4976 \$5097 \$5837 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1957 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1958 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1959 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1960 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1961 \$5838 \$5853 \$5833 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1962 \$5100 \$5853 \$5838 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1963 \$5839 \$5853 \$5186 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1964 \$5840 \$5853 \$5839 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1965 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1966 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1967 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1968 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1969 \$5841 \$5119 \$5120 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1970 \$2147 \$5119 \$5841 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1971 \$5842 \$5958 \$2147 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1972 \$5853 \$5958 \$5842 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1973 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1974 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1975 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1976 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1977 \$5843 \$5105 \$5105 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1978 VDD \$5105 \$5843 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1979 \$5844 \$5105 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1980 \$4977 \$5105 \$5844 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1981 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1982 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1983 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1984 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1985 \$5845 \$5854 \$5840 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1986 \$5108 \$5854 \$5845 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1987 \$5846 \$5854 \$5187 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1988 B1 \$5854 \$5846 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1989 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1990 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1991 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1992 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1993 \$5848 \$5121 \$5122 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1994 \$2150 \$5121 \$5848 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1995 \$5849 \$5959 \$2150 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1996 \$5854 \$5959 \$5849 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1997 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1998 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1999 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2000 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2001 \$5975 \$5073 \$4973 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2002 VDD \$5073 \$5975 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2003 \$5976 \$5073 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2004 \$5073 \$5073 \$5976 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2005 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2006 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2007 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2008 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2009 \$5977 \$5850 \$5955 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2010 VSS \$5850 \$5977 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2011 \$5978 \$5850 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2012 \$5955 \$5850 \$5978 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2013 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2014 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2015 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2016 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2017 \$5979 \$5955 \$5850 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2018 \$3943 \$5955 \$5979 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2019 \$5980 \$5113 \$3943 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2020 \$5114 \$5113 \$5980 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2021 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2022 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2023 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2024 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2025 \$5981 \$5081 \$4974 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2026 VDD \$5081 \$5981 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2027 \$5982 \$5081 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2028 \$5081 \$5081 \$5982 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2029 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2030 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2031 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2032 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2033 \$5983 \$5851 \$5956 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2034 VSS \$5851 \$5983 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2035 \$5984 \$5851 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2036 \$5956 \$5851 \$5984 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2037 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2038 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2039 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2040 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2041 \$5985 \$5956 \$5851 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2042 \$3944 \$5956 \$5985 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2043 \$5986 \$5115 \$3944 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2044 \$5116 \$5115 \$5986 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2045 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2046 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2047 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2048 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2049 \$5987 \$5089 \$4975 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2050 VDD \$5089 \$5987 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2051 \$5988 \$5089 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2052 \$5089 \$5089 \$5988 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2053 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2054 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2055 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2056 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2057 \$5989 \$5852 \$5957 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2058 VSS \$5852 \$5989 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2059 \$5990 \$5852 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2060 \$5957 \$5852 \$5990 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2061 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2062 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2063 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2064 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2065 \$5991 \$5957 \$5852 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2066 \$3945 \$5957 \$5991 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2067 \$5992 \$5117 \$3945 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2068 \$5118 \$5117 \$5992 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2069 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2070 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2071 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2072 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2073 \$5993 \$5097 \$4976 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2074 VDD \$5097 \$5993 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2075 \$5994 \$5097 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2076 \$5097 \$5097 \$5994 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2077 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2078 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2079 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2080 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2081 \$5995 \$5853 \$5958 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2082 VSS \$5853 \$5995 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2083 \$5996 \$5853 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2084 \$5958 \$5853 \$5996 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2085 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2086 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2087 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2088 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2089 \$5997 \$5958 \$5853 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2090 \$2147 \$5958 \$5997 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2091 \$5998 \$5119 \$2147 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2092 \$5120 \$5119 \$5998 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2093 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2094 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2095 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2096 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2097 \$5999 \$5105 \$4977 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2098 VDD \$5105 \$5999 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2099 \$6000 \$5105 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2100 \$5105 \$5105 \$6000 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2101 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2102 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2103 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2104 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2105 \$6001 \$5854 \$5959 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2106 VSS \$5854 \$6001 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2107 \$6002 \$5854 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2108 \$5959 \$5854 \$6002 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2109 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2110 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2111 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2112 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2113 \$6003 \$5959 \$5854 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2114 \$2150 \$5959 \$6003 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2115 \$6004 \$5121 \$2150 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2116 \$5122 \$5121 \$6004 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2117 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2118 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2119 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2120 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2121 \$6110 \$5073 \$5073 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2122 VDD \$5073 \$6110 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2123 \$6111 \$5073 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2124 \$4973 \$5073 \$6111 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2125 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2126 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2127 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2128 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2129 \$6112 \$5850 \$5955 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2130 VSS \$5850 \$6112 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2131 \$6113 \$5850 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2132 \$5955 \$5850 \$6113 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2133 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2134 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2135 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2136 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2137 \$6114 \$5113 \$5114 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2138 \$3943 \$5113 \$6114 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2139 \$6115 \$5955 \$3943 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2140 \$5850 \$5955 \$6115 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2141 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2142 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2143 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2144 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2145 \$6116 \$5081 \$5081 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2146 VDD \$5081 \$6116 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2147 \$6117 \$5081 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2148 \$4974 \$5081 \$6117 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2149 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2150 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2151 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2152 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2153 \$6118 \$5851 \$5956 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2154 VSS \$5851 \$6118 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2155 \$6119 \$5851 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2156 \$5956 \$5851 \$6119 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2157 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2158 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2159 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2160 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2161 \$6120 \$5115 \$5116 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2162 \$3944 \$5115 \$6120 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2163 \$6121 \$5956 \$3944 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2164 \$5851 \$5956 \$6121 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2165 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2166 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2167 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2168 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2169 \$6122 \$5089 \$5089 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2170 VDD \$5089 \$6122 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2171 \$6123 \$5089 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2172 \$4975 \$5089 \$6123 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2173 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2174 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2175 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2176 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2177 \$6124 \$5852 \$5957 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2178 VSS \$5852 \$6124 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2179 \$6125 \$5852 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2180 \$5957 \$5852 \$6125 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2181 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2182 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2183 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2184 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2185 \$6126 \$5117 \$5118 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2186 \$3945 \$5117 \$6126 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2187 \$6127 \$5957 \$3945 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2188 \$5852 \$5957 \$6127 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2189 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2190 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2191 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2192 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2193 \$6128 \$5097 \$5097 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2194 VDD \$5097 \$6128 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2195 \$6129 \$5097 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2196 \$4976 \$5097 \$6129 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2197 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2198 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2199 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2200 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2201 \$6130 \$5853 \$5958 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2202 VSS \$5853 \$6130 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2203 \$6131 \$5853 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2204 \$5958 \$5853 \$6131 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2205 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2206 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2207 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2208 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2209 \$6132 \$5119 \$5120 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2210 \$2147 \$5119 \$6132 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2211 \$6133 \$5958 \$2147 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2212 \$5853 \$5958 \$6133 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2213 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2214 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2215 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2216 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2217 \$6134 \$5105 \$5105 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2218 VDD \$5105 \$6134 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2219 \$6135 \$5105 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2220 \$4977 \$5105 \$6135 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2221 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2222 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2223 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2224 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2225 \$6136 \$5854 \$5959 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2226 VSS \$5854 \$6136 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2227 \$6137 \$5854 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2228 \$5959 \$5854 \$6137 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2229 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2230 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2231 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2232 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2233 \$6138 \$5121 \$5122 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2234 \$2150 \$5121 \$6138 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2235 \$6139 \$5959 \$2150 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2236 \$5854 \$5959 \$6139 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2237 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2238 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2239 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2240 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2241 \$6270 \$5073 \$4973 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2242 VDD \$5073 \$6270 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2243 \$6271 \$5073 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2244 \$5073 \$5073 \$6271 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2245 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2246 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2247 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2248 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2249 \$6272 \$5850 \$5819 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2250 \$5183 \$5850 \$6272 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2251 \$6273 \$5850 \$5076 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2252 A1 \$5850 \$6273 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2253 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2254 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2255 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2256 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2257 \$6274 \$5955 \$5850 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2258 \$3943 \$5955 \$6274 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2259 \$6275 \$5113 \$3943 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2260 \$5114 \$5113 \$6275 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2261 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2262 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2263 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2264 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2265 \$6276 \$5081 \$4974 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2266 VDD \$5081 \$6276 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2267 \$6277 \$5081 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2268 \$5081 \$5081 \$6277 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2269 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2270 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2271 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2272 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2273 \$6278 \$5851 \$5826 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2274 \$5184 \$5851 \$6278 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2275 \$6279 \$5851 \$5084 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2276 \$5819 \$5851 \$6279 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2277 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2278 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2279 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2280 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2281 \$6280 \$5956 \$5851 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2282 \$3944 \$5956 \$6280 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2283 \$6281 \$5115 \$3944 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2284 \$5116 \$5115 \$6281 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2285 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2286 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2287 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2288 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2289 \$6282 \$5089 \$4975 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2290 VDD \$5089 \$6282 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2291 \$6283 \$5089 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2292 \$5089 \$5089 \$6283 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2293 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2294 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2295 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2296 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2297 \$6284 \$5852 \$5833 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2298 \$5185 \$5852 \$6284 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2299 \$6285 \$5852 \$5092 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2300 \$5826 \$5852 \$6285 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2301 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2302 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2303 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2304 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2305 \$6286 \$5957 \$5852 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2306 \$3945 \$5957 \$6286 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2307 \$6287 \$5117 \$3945 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2308 \$5118 \$5117 \$6287 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2309 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2310 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2311 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2312 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2313 \$6288 \$5097 \$4976 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2314 VDD \$5097 \$6288 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2315 \$6289 \$5097 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2316 \$5097 \$5097 \$6289 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2317 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2318 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2319 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2320 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2321 \$6290 \$5853 \$5840 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2322 \$5186 \$5853 \$6290 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2323 \$6291 \$5853 \$5100 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2324 \$5833 \$5853 \$6291 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2325 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2326 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2327 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2328 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2329 \$6292 \$5958 \$5853 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2330 \$2147 \$5958 \$6292 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2331 \$6293 \$5119 \$2147 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2332 \$5120 \$5119 \$6293 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2333 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2334 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2335 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2336 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2337 \$6294 \$5105 \$4977 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2338 VDD \$5105 \$6294 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2339 \$6295 \$5105 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2340 \$5105 \$5105 \$6295 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2341 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2342 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2343 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2344 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2345 \$6296 \$5854 B1 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2346 \$5187 \$5854 \$6296 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2347 \$6297 \$5854 \$5108 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2348 \$5840 \$5854 \$6297 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2349 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2350 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2351 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2352 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2353 \$6298 \$5959 \$5854 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2354 \$2150 \$5959 \$6298 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2355 \$6299 \$5121 \$2150 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2356 \$5122 \$5121 \$6299 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2357 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2358 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2359 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2360 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2361 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2362 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2363 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2364 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2365 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2366 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2367 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2368 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2369 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2370 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2371 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2372 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2373 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2374 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2375 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2376 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2377 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2378 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2379 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2380 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2381 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2382 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2383 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2384 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2385 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2386 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2387 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2388 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2389 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2390 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2391 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2392 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2393 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2394 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2395 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2396 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2397 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2398 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2399 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2400 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2401 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2402 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2403 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2404 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2405 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2406 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2407 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2408 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2409 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2410 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2411 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2412 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2413 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2414 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2415 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2416 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2417 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2418 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2419 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2420 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2421 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2422 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2423 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2424 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2425 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2426 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2427 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2428 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2429 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2430 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2431 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2432 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2433 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2434 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2435 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2436 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2437 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2438 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2439 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2440 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2441 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2442 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2443 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2444 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2445 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2446 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2447 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2448 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2449 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2450 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2451 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2452 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2453 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2454 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2455 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2456 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2457 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2458 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2459 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2460 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2461 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2462 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2463 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2464 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2465 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2466 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2467 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2468 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2469 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2470 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2471 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2472 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2473 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2474 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2475 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2476 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2477 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2478 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2479 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2480 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2481 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2482 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2483 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2484 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2485 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2486 AVDD IREF \$9382 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2487 \$9382 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2488 AVDD IREF \$9382 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2489 \$9382 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2490 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2491 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2492 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2493 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2494 AVDD IREF \$8587 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2495 \$8587 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2496 AVDD IREF \$8587 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2497 \$8587 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2498 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2499 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2500 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2501 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2502 AVDD IREF \$8587 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2503 \$8587 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2504 AVDD IREF \$8587 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2505 \$8587 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2506 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2507 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2508 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2509 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2510 AVDD IREF \$9382 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2511 \$9382 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2512 AVDD IREF \$9382 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2513 \$9382 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2514 AVDD IREF \$8587 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2515 \$8587 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2516 AVDD IREF \$8587 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2517 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2518 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2519 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2520 \$9382 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2521 AVDD IREF \$9382 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2522 \$9382 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2523 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2524 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2525 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2526 AVDD IREF \$9382 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2527 \$9382 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2528 AVDD IREF \$9382 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2529 \$8587 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2530 AVDD IREF \$8587 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2531 \$8587 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2532 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2533 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2534 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2535 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2536 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2537 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2538 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2539 AVDD IREF \$9382 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2540 \$9382 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2541 AVDD IREF \$9382 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2542 \$9382 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2543 AVDD IREF \$8587 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2544 \$8587 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2545 AVDD IREF \$8587 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2546 \$8587 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2547 AVDD IREF \$9382 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2548 \$9382 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2549 AVDD IREF \$9382 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2550 \$9382 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2551 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2552 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2553 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2554 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2555 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2556 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2557 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2558 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2559 AVDD IREF \$8587 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2560 \$8587 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2561 AVDD IREF \$8587 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2562 \$8587 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2563 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2564 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2565 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2566 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2567 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2568 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2569 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2570 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2571 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2572 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2573 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2574 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2575 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2576 \$14597 \$8078 \$13791 AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P
+ PS=3.7U PD=2.04U
M$2577 \$14598 \$8078 \$14597 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P
+ PS=2.04U PD=2.04U
M$2578 \$14599 \$8078 \$14598 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P
+ PS=2.04U PD=3.7U
M$2579 \$12709 \$8078 \$12708 AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P
+ PS=3.7U PD=2.04U
M$2580 \$12710 \$8078 \$12709 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P
+ PS=2.04U PD=2.04U
M$2581 AVDD \$8078 \$12710 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P
+ PS=2.04U PD=3.7U
M$2582 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P PS=3.7U
+ PD=2.04U
M$2583 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P PS=2.04U
+ PD=2.04U
M$2584 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P PS=2.04U
+ PD=3.7U
M$2585 \$13385 \$8078 \$12708 AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P
+ PS=3.7U PD=2.04U
M$2586 \$13386 \$8078 \$13385 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P
+ PS=2.04U PD=2.04U
M$2587 \$13387 \$8078 \$13386 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P
+ PS=2.04U PD=3.7U
M$2588 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P PS=3.7U
+ PD=2.04U
M$2589 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P PS=2.04U
+ PD=2.04U
M$2590 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P PS=2.04U
+ PD=3.7U
M$2591 \$13792 \$8078 \$13791 AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P
+ PS=3.7U PD=2.04U
M$2592 \$13793 \$8078 \$13792 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P
+ PS=2.04U PD=2.04U
M$2593 \$13387 \$8078 \$13793 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P
+ PS=2.04U PD=3.7U
M$2594 \$8078 \$8078 \$14599 AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P
+ PS=3.7U PD=3.7U
M$2595 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2596 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2597 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2598 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2599 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2600 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2601 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2602 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2603 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2604 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2605 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$2606 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2607 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2608 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2609 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2610 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2611 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2612 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2613 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2614 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2615 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2616 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2617 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2618 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2619 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2620 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2621 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2622 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2623 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2624 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2625 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2626 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2627 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2628 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2629 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2630 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2631 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2632 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2633 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2634 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2635 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2636 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2637 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2638 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2639 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2640 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2641 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2642 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2643 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2644 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2645 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2646 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2647 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2648 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2649 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2650 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2651 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2652 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2653 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2654 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2655 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2656 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2657 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2658 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2659 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2660 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2661 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2662 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2663 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2664 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2665 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2666 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2667 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2668 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2669 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2670 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2671 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2672 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2673 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2674 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2675 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2676 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2677 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2678 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2679 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2680 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2681 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2682 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2683 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2684 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2685 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2686 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2687 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2688 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2689 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2690 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2691 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2692 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2693 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2694 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2695 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2696 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2697 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2698 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2699 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2700 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2701 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2702 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2703 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2704 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2705 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2706 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2707 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2708 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2709 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2710 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2711 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2712 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2713 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2714 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2715 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2716 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2717 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2718 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2719 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2720 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2721 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2722 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2723 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2724 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2725 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2726 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2727 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2728 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2729 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2730 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2731 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2732 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2733 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2734 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2735 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2736 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2737 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2738 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2739 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2740 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2741 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2742 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2743 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2744 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2745 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2746 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2747 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2748 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2749 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2750 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2751 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2752 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2753 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2754 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2755 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2756 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2757 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2758 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2759 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2760 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2761 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2762 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2763 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2764 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2765 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2766 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2767 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2768 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2769 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2770 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2771 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2772 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2773 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2774 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2775 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2776 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2777 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2778 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2779 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2780 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2781 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2782 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2783 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2784 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2785 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2786 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2787 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2788 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2789 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2790 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2791 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2792 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2793 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2794 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2795 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2796 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2797 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2798 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2799 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2800 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2801 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2802 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2803 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2804 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2805 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2806 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2807 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2808 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2809 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2810 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2811 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2812 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2813 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2814 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2815 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2816 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2817 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2818 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2819 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2820 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2821 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2822 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2823 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2824 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2825 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2826 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2827 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2828 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2829 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2830 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2831 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2832 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2833 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2834 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2835 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2836 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2837 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2838 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2839 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2840 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2841 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2842 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2843 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2844 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2845 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2846 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2847 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2848 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2849 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2850 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2851 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2852 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2853 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2854 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2855 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2856 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2857 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2858 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2859 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2860 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2861 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2862 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2863 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2864 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2865 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2866 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2867 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2868 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2869 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2870 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2871 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2872 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2873 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2874 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2875 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2876 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$2877 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$2878 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2879 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2880 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2881 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2882 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2883 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2884 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2885 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2886 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2887 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2888 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2889 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2890 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2891 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2892 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2893 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2894 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2895 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2896 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2897 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2898 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2899 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2900 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2901 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2902 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2903 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2904 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2905 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2906 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2907 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2908 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2909 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2910 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2911 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2912 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2913 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2914 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2915 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2916 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2917 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2918 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2919 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2920 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2921 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2922 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2923 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2924 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2925 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2926 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2927 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2928 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2929 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2930 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2931 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2932 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2933 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2934 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2935 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2936 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2937 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2938 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2939 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2940 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2941 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2942 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2943 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2944 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2945 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2946 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2947 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2948 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2949 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2950 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2951 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2952 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2953 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2954 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2955 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2956 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2957 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2958 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2959 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2960 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2961 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2962 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2963 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2964 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2965 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2966 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2967 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2968 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2969 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2970 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2971 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2972 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2973 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2974 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2975 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2976 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2977 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2978 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2979 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2980 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2981 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$2982 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2983 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2984 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2985 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2986 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2987 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2988 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2989 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2990 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2991 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2992 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2993 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2994 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$2995 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2996 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2997 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$2998 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$2999 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3000 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3001 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3002 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3003 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3004 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3005 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3006 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3007 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3008 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3009 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3010 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3011 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3012 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3013 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3014 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3015 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3016 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3017 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3018 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3019 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3020 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3021 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3022 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3023 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3024 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3025 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3026 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3027 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3028 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3029 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3030 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3031 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3032 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3033 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3034 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3035 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3036 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3037 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3038 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3039 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3040 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3041 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3042 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3043 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3044 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3045 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3046 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3047 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3048 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3049 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3050 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3051 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3052 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3053 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3054 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3055 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3056 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3057 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3058 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3059 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3060 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3061 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3062 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3063 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3064 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3065 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3066 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3067 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3068 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3069 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3070 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3071 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3072 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3073 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3074 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3075 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3076 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3077 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3078 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3079 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3080 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3081 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3082 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3083 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3084 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3085 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3086 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3087 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3088 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3089 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3090 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3091 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3092 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3093 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3094 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3095 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3096 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3097 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3098 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3099 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3100 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3101 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3102 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3103 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3104 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3105 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3106 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3107 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3108 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3109 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3110 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3111 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3112 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3113 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3114 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3115 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3116 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3117 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3118 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3119 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3120 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3121 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3122 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3123 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3124 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3125 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3126 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3127 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3128 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3129 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3130 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3131 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3132 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3133 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3134 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3135 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3136 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3137 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3138 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3139 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3140 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3141 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3142 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3143 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3144 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3145 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3146 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3147 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3148 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3149 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3150 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3151 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3152 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3153 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3154 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3155 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3156 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3157 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3158 \$22196 VN \$7408 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3159 \$7408 VN \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3160 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3161 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3162 \$22196 VP \$7673 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3163 \$7673 VP \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3164 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3165 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3166 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3167 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3168 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3169 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3170 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3171 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3172 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3173 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3174 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3175 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3176 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3177 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3178 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3179 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3180 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3181 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3182 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3183 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3184 \$22198 \$8078 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3185 VOUT \$8078 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3186 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3187 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3188 \$22197 \$8078 \$14873 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P
+ PS=2.84U PD=2.84U
M$3189 \$14873 \$8078 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P
+ PS=2.84U PD=5.3U
M$3190 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3191 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3192 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3193 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3194 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3195 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3196 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3197 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3198 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3199 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3200 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3201 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3202 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3203 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3204 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3205 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3206 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3207 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3208 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3209 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3210 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3211 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3212 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3213 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3214 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3215 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3216 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3217 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3218 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3219 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3220 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3221 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3222 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3223 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3224 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3225 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3226 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3227 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3228 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3229 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3230 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3231 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3232 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3233 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3234 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3235 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3236 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3237 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3238 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3239 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3240 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3241 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3242 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3243 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3244 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3245 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3246 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3247 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3248 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3249 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3250 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3251 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3252 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3253 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3254 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3255 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3256 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3257 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3258 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3259 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3260 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3261 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3262 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3263 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3264 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3265 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3266 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3267 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3268 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3269 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3270 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3271 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3272 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3273 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3274 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3275 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3276 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3277 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3278 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3279 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3280 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3281 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3282 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3283 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3284 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3285 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3286 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3287 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3288 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3289 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3290 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3291 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3292 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3293 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3294 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3295 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3296 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3297 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3298 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3299 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3300 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3301 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3302 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3303 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3304 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3305 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3306 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3307 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3308 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3309 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3310 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3311 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3312 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3313 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3314 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3315 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3316 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3317 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3318 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3319 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3320 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3321 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3322 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3323 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3324 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3325 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3326 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3327 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3328 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3329 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3330 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3331 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3332 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3333 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3334 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3335 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3336 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3337 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3338 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3339 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3340 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3341 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3342 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3343 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3344 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3345 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3346 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3347 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3348 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3349 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3350 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3351 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3352 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3353 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3354 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3355 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3356 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3357 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3358 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3359 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3360 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3361 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3362 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3363 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3364 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3365 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3366 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3367 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3368 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3369 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3370 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3371 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3372 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3373 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3374 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3375 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3376 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3377 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3378 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3379 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3380 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3381 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3382 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3383 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3384 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3385 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3386 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3387 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3388 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3389 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3390 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3391 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3392 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3393 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3394 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3395 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3396 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3397 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3398 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3399 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3400 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3401 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3402 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3403 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3404 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3405 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3406 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3407 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3408 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3409 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3410 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3411 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3412 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3413 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3414 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3415 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3416 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3417 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3418 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3419 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3420 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3421 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3422 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3423 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3424 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3425 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3426 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3427 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3428 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3429 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3430 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3431 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3432 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3433 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3434 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3435 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3436 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3437 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3438 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3439 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3440 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3441 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3442 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3443 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3444 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3445 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3446 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3447 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3448 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3449 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3450 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3451 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3452 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3453 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3454 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3455 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3456 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3457 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3458 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3459 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3460 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3461 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3462 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3463 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3464 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3465 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3466 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3467 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3468 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3469 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3470 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3471 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3472 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3473 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3474 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3475 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3476 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3477 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3478 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3479 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3480 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3481 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3482 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3483 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3484 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3485 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3486 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3487 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3488 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3489 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3490 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3491 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3492 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3493 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3494 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3495 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3496 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3497 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3498 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3499 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3500 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3501 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3502 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3503 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3504 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3505 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3506 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3507 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3508 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3509 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3510 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3511 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3512 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3513 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3514 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3515 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3516 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3517 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3518 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3519 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3520 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3521 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3522 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3523 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3524 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3525 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3526 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3527 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3528 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3529 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3530 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3531 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3532 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3533 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3534 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3535 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3536 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3537 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3538 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3539 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3540 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3541 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3542 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3543 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3544 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3545 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3546 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3547 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3548 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3549 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3550 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3551 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3552 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3553 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3554 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3555 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3556 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3557 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3558 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3559 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3560 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3561 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3562 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3563 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3564 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3565 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3566 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3567 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3568 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3569 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3570 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3571 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3572 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3573 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3574 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3575 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3576 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3577 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3578 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3579 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3580 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3581 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3582 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3583 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3584 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3585 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3586 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3587 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3588 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3589 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3590 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3591 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3592 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3593 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3594 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3595 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3596 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3597 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3598 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3599 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3600 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3601 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3602 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3603 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3604 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3605 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3606 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3607 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3608 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3609 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3610 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3611 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3612 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3613 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3614 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3615 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3616 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3617 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3618 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3619 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3620 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3621 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3622 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3623 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3624 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3625 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3626 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3627 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3628 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3629 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3630 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3631 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3632 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3633 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3634 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3635 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3636 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3637 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3638 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3639 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3640 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3641 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3642 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3643 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3644 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3645 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3646 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3647 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3648 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3649 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3650 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3651 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3652 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3653 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3654 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3655 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3656 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3657 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3658 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3659 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3660 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3661 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3662 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3663 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3664 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3665 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3666 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3667 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3668 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3669 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3670 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3671 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3672 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3673 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3674 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3675 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3676 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3677 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3678 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3679 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3680 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3681 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3682 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3683 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3684 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3685 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3686 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3687 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3688 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3689 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3690 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3691 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3692 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3693 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3694 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3695 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3696 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3697 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3698 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3699 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3700 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3701 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3702 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3703 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3704 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3705 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3706 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3707 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3708 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3709 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3710 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3711 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3712 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3713 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3714 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3715 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3716 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3717 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3718 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3719 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3720 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3721 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3722 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3723 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3724 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3725 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3726 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3727 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3728 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3729 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3730 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3731 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3732 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3733 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3734 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3735 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3736 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3737 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3738 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3739 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3740 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3741 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3742 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3743 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3744 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3745 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3746 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3747 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3748 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3749 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3750 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3751 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3752 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3753 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3754 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3755 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3756 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3757 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3758 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3759 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3760 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3761 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3762 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3763 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3764 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3765 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3766 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3767 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3768 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3769 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3770 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3771 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3772 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3773 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3774 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3775 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3776 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3777 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3778 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3779 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3780 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3781 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3782 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3783 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3784 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3785 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3786 AVDD IREF \$22196 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3787 \$22196 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3788 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3789 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3790 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3791 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3792 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3793 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3794 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3795 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3796 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3797 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3798 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3799 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3800 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3801 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3802 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3803 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3804 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3805 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3806 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3807 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3808 AVDD \$14873 \$22198 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3809 \$22198 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3810 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$3811 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3812 AVDD \$14873 \$22197 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3813 \$22197 \$14873 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$3814 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3815 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3816 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3817 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3818 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3819 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3820 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3821 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3822 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3823 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3824 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3825 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3826 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3827 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3828 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3829 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3830 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3831 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3832 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3833 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3834 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3835 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3836 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3837 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3838 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3839 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3840 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3841 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3842 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3843 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3844 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3845 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3846 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3847 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3848 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3849 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3850 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3851 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3852 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3853 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3854 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3855 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3856 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3857 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3858 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3859 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3860 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3861 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3862 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3863 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3864 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$3865 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3866 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$3867 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3868 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3869 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3870 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3871 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3872 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3873 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3874 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3875 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3876 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3877 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3878 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3879 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3880 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3881 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3882 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3883 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3884 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3885 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3886 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3887 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3888 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3889 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3890 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3891 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3892 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3893 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3894 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3895 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3896 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3897 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3898 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3899 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3900 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3901 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3902 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3903 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3904 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3905 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3906 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3907 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3908 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3909 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3910 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3911 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3912 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3913 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3914 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3915 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3916 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3917 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3918 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3919 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3920 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3921 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3922 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3923 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3924 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3925 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3926 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3927 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3928 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3929 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3930 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3931 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3932 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3933 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3934 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3935 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3936 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3937 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3938 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3939 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3940 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3941 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3942 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3943 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3944 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3945 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3946 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3947 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3948 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3949 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3950 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3951 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3952 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3953 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3954 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3955 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3956 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3957 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3958 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3959 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3960 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3961 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3962 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3963 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3964 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3965 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3966 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3967 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3968 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3969 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3970 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3971 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3972 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3973 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3974 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3975 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3976 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3977 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3978 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3979 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3980 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3981 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3982 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3983 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3984 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3985 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3986 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3987 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3988 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3989 \$886 \$916 \$917 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$3990 \$866 \$916 \$886 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$3991 \$887 \$259 \$866 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$3992 \$173 \$259 \$887 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$3993 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3994 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3995 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3996 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$3997 \$888 \$917 \$139 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$3998 \$259 \$917 \$888 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$3999 \$889 \$917 \$259 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4000 \$116 \$917 \$889 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4001 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4002 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4003 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4004 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4005 \$890 \$258 \$25 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4006 VSS \$258 \$890 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4007 \$891 \$258 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4008 \$258 \$258 \$891 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4009 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4010 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4011 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4012 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4013 \$892 \$918 \$919 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4014 \$867 \$918 \$892 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4015 \$893 \$261 \$867 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4016 \$175 \$261 \$893 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4017 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4018 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4019 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4020 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4021 \$894 \$919 \$147 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4022 \$261 \$919 \$894 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4023 \$895 \$919 \$261 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4024 \$117 \$919 \$895 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4025 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4026 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4027 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4028 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4029 \$896 \$260 \$26 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4030 VSS \$260 \$896 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4031 \$897 \$260 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4032 \$260 \$260 \$897 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4033 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4034 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4035 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4036 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4037 \$898 \$920 \$921 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4038 \$868 \$920 \$898 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4039 \$899 \$263 \$868 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4040 \$177 \$263 \$899 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4041 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4042 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4043 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4044 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4045 \$900 \$921 \$154 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4046 \$263 \$921 \$900 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4047 \$901 \$921 \$263 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4048 \$118 \$921 \$901 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4049 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4050 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4051 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4052 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4053 \$902 \$262 \$27 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4054 VSS \$262 \$902 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4055 \$903 \$262 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4056 \$262 \$262 \$903 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4057 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4058 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4059 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4060 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4061 \$904 \$922 \$923 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4062 \$869 \$922 \$904 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4063 \$905 \$265 \$869 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4064 \$179 \$265 \$905 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4065 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4066 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4067 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4068 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4069 \$906 \$923 \$161 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4070 \$265 \$923 \$906 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4071 \$907 \$923 \$265 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4072 \$119 \$923 \$907 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4073 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4074 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4075 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4076 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4077 \$908 \$264 \$28 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4078 VSS \$264 \$908 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4079 \$909 \$264 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4080 \$264 \$264 \$909 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4081 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4082 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4083 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4084 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4085 \$910 \$924 \$925 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4086 \$870 \$924 \$910 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4087 \$911 \$267 \$870 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4088 \$181 \$267 \$911 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4089 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4090 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4091 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4092 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4093 \$912 \$925 \$169 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4094 \$267 \$925 \$912 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4095 \$913 \$925 \$267 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4096 \$120 \$925 \$913 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4097 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4098 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4099 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4100 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4101 \$914 \$266 \$29 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4102 VSS \$266 \$914 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4103 \$915 \$266 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4104 \$266 \$266 \$915 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4105 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4106 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4107 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4108 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4109 \$1041 \$259 \$173 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4110 \$866 \$259 \$1041 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4111 \$1042 \$916 \$866 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4112 \$917 \$916 \$1042 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4113 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4114 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4115 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4116 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4117 \$1043 \$917 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4118 \$916 \$917 \$1043 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4119 \$1044 \$917 \$916 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4120 VDD \$917 \$1044 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4121 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4122 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4123 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4124 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4125 \$1045 \$258 \$258 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4126 VSS \$258 \$1045 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4127 \$1046 \$258 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4128 \$25 \$258 \$1046 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4129 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4130 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4131 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4132 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4133 \$1047 \$261 \$175 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4134 \$867 \$261 \$1047 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4135 \$1048 \$918 \$867 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4136 \$919 \$918 \$1048 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4137 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4138 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4139 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4140 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4141 \$1049 \$919 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4142 \$918 \$919 \$1049 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4143 \$1050 \$919 \$918 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4144 VDD \$919 \$1050 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4145 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4146 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4147 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4148 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4149 \$1051 \$260 \$260 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4150 VSS \$260 \$1051 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4151 \$1052 \$260 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4152 \$26 \$260 \$1052 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4153 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4154 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4155 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4156 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4157 \$1053 \$263 \$177 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4158 \$868 \$263 \$1053 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4159 \$1054 \$920 \$868 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4160 \$921 \$920 \$1054 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4161 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4162 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4163 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4164 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4165 \$1055 \$921 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4166 \$920 \$921 \$1055 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4167 \$1056 \$921 \$920 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4168 VDD \$921 \$1056 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4169 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4170 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4171 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4172 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4173 \$1057 \$262 \$262 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4174 VSS \$262 \$1057 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4175 \$1058 \$262 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4176 \$27 \$262 \$1058 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4177 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4178 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4179 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4180 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4181 \$1059 \$265 \$179 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4182 \$869 \$265 \$1059 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4183 \$1060 \$922 \$869 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4184 \$923 \$922 \$1060 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4185 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4186 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4187 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4188 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4189 \$1061 \$923 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4190 \$922 \$923 \$1061 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4191 \$1062 \$923 \$922 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4192 VDD \$923 \$1062 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4193 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4194 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4195 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4196 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4197 \$1063 \$264 \$264 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4198 VSS \$264 \$1063 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4199 \$1064 \$264 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4200 \$28 \$264 \$1064 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4201 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4202 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4203 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4204 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4205 \$1065 \$267 \$181 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4206 \$870 \$267 \$1065 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4207 \$1066 \$924 \$870 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4208 \$925 \$924 \$1066 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4209 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4210 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4211 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4212 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4213 \$1067 \$925 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4214 \$924 \$925 \$1067 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4215 \$1068 \$925 \$924 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4216 VDD \$925 \$1068 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4217 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4218 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4219 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4220 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4221 \$1069 \$266 \$266 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4222 VSS \$266 \$1069 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4223 \$1070 \$266 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4224 \$29 \$266 \$1070 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4225 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4226 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4227 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4228 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4229 \$1176 \$916 \$917 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4230 \$866 \$916 \$1176 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4231 \$1177 \$259 \$866 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4232 \$173 \$259 \$1177 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4233 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4234 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4235 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4236 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4237 \$1178 \$917 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4238 \$916 \$917 \$1178 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4239 \$1179 \$917 \$916 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4240 VDD \$917 \$1179 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4241 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4242 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4243 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4244 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4245 \$1180 \$258 \$25 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4246 VSS \$258 \$1180 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4247 \$1181 \$258 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4248 \$258 \$258 \$1181 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4249 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4250 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4251 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4252 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4253 \$1182 \$918 \$919 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4254 \$867 \$918 \$1182 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4255 \$1183 \$261 \$867 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4256 \$175 \$261 \$1183 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4257 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4258 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4259 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4260 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4261 \$1184 \$919 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4262 \$918 \$919 \$1184 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4263 \$1185 \$919 \$918 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4264 VDD \$919 \$1185 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4265 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4266 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4267 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4268 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4269 \$1186 \$260 \$26 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4270 VSS \$260 \$1186 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4271 \$1187 \$260 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4272 \$260 \$260 \$1187 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4273 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4274 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4275 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4276 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4277 \$1188 \$920 \$921 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4278 \$868 \$920 \$1188 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4279 \$1189 \$263 \$868 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4280 \$177 \$263 \$1189 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4281 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4282 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4283 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4284 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4285 \$1190 \$921 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4286 \$920 \$921 \$1190 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4287 \$1191 \$921 \$920 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4288 VDD \$921 \$1191 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4289 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4290 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4291 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4292 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4293 \$1192 \$262 \$27 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4294 VSS \$262 \$1192 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4295 \$1193 \$262 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4296 \$262 \$262 \$1193 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4297 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4298 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4299 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4300 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4301 \$1194 \$922 \$923 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4302 \$869 \$922 \$1194 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4303 \$1195 \$265 \$869 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4304 \$179 \$265 \$1195 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4305 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4306 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4307 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4308 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4309 \$1196 \$923 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4310 \$922 \$923 \$1196 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4311 \$1197 \$923 \$922 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4312 VDD \$923 \$1197 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4313 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4314 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4315 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4316 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4317 \$1198 \$264 \$28 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4318 VSS \$264 \$1198 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4319 \$1199 \$264 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4320 \$264 \$264 \$1199 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4321 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4322 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4323 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4324 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4325 \$1200 \$924 \$925 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4326 \$870 \$924 \$1200 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4327 \$1201 \$267 \$870 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4328 \$181 \$267 \$1201 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4329 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4330 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4331 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4332 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4333 \$1202 \$925 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4334 \$924 \$925 \$1202 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4335 \$1203 \$925 \$924 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4336 VDD \$925 \$1203 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4337 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4338 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4339 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4340 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4341 \$1204 \$266 \$29 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4342 VSS \$266 \$1204 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4343 \$1205 \$266 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4344 \$266 \$266 \$1205 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4345 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4346 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4347 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4348 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4349 \$1321 \$259 \$173 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4350 \$866 \$259 \$1321 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4351 \$1322 \$916 \$866 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4352 \$917 \$916 \$1322 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4353 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4354 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4355 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4356 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4357 \$1323 \$917 \$116 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4358 \$259 \$917 \$1323 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4359 \$1324 \$917 \$259 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4360 \$139 \$917 \$1324 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4361 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4362 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4363 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4364 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4365 \$1325 \$258 \$258 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4366 VSS \$258 \$1325 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4367 \$1326 \$258 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4368 \$25 \$258 \$1326 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4369 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4370 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4371 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4372 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4373 \$1327 \$261 \$175 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4374 \$867 \$261 \$1327 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4375 \$1328 \$918 \$867 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4376 \$919 \$918 \$1328 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4377 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4378 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4379 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4380 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4381 \$1329 \$919 \$117 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4382 \$261 \$919 \$1329 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4383 \$1330 \$919 \$261 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4384 \$147 \$919 \$1330 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4385 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4386 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4387 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4388 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4389 \$1331 \$260 \$260 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4390 VSS \$260 \$1331 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4391 \$1332 \$260 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4392 \$26 \$260 \$1332 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4393 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4394 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4395 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4396 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4397 \$1333 \$263 \$177 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4398 \$868 \$263 \$1333 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4399 \$1334 \$920 \$868 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4400 \$921 \$920 \$1334 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4401 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4402 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4403 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4404 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4405 \$1335 \$921 \$118 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4406 \$263 \$921 \$1335 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4407 \$1336 \$921 \$263 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4408 \$154 \$921 \$1336 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4409 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4410 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4411 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4412 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4413 \$1337 \$262 \$262 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4414 VSS \$262 \$1337 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4415 \$1338 \$262 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4416 \$27 \$262 \$1338 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4417 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4418 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4419 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4420 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4421 \$1339 \$265 \$179 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4422 \$869 \$265 \$1339 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4423 \$1340 \$922 \$869 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4424 \$923 \$922 \$1340 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4425 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4426 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4427 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4428 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4429 \$1341 \$923 \$119 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4430 \$265 \$923 \$1341 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4431 \$1342 \$923 \$265 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4432 \$161 \$923 \$1342 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4433 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4434 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4435 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4436 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4437 \$1343 \$264 \$264 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4438 VSS \$264 \$1343 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4439 \$1344 \$264 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4440 \$28 \$264 \$1344 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4441 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4442 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4443 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4444 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4445 \$1345 \$267 \$181 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4446 \$870 \$267 \$1345 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4447 \$1346 \$924 \$870 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4448 \$925 \$924 \$1346 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4449 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4450 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4451 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4452 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4453 \$1347 \$925 \$120 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4454 \$267 \$925 \$1347 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4455 \$1348 \$925 \$267 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4456 \$169 \$925 \$1348 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4457 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4458 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4459 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4460 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4461 \$1349 \$266 \$266 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4462 VSS \$266 \$1349 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4463 \$1350 \$266 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4464 \$29 \$266 \$1350 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4465 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4466 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4467 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4468 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4469 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4470 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4471 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4472 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4473 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4474 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4475 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4476 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4477 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4478 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4479 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4480 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4481 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4482 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4483 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4484 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4485 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4486 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4487 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4488 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4489 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4490 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4491 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4492 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4493 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4494 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4495 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4496 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4497 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4498 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4499 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4500 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4501 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4502 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4503 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4504 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4505 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4506 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4507 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4508 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4509 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4510 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4511 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4512 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4513 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4514 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4515 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4516 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4517 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4518 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4519 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4520 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4521 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4522 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4523 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4524 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4525 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4526 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4527 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4528 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4529 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4530 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4531 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4532 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4533 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4534 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4535 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4536 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4537 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4538 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4539 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4540 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4541 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4542 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4543 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4544 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4545 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4546 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4547 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4548 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4549 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4550 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4551 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4552 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4553 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4554 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4555 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4556 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4557 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4558 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4559 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4560 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4561 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4562 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4563 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4564 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4565 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4566 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4567 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4568 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4569 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4570 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4571 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4572 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4573 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4574 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4575 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4576 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4577 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4578 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4579 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4580 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4581 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4582 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4583 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4584 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4585 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4586 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4587 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4588 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4589 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4590 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4591 \$1781 \$1773 \$1780 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4592 \$916 \$1773 \$1781 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4593 \$1783 \$1773 \$1782 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4594 \$1784 \$1773 \$1783 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4595 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4596 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4597 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4598 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4599 \$1785 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4600 \$1786 \$1773 \$1785 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4601 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4602 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4603 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4604 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4605 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4606 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4607 \$1788 \$1773 \$1787 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4608 \$918 \$1773 \$1788 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4609 \$1790 \$1773 \$1789 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4610 \$1791 \$1773 \$1790 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4611 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4612 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4613 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4614 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4615 \$1792 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4616 \$1793 \$1773 \$1792 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4617 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4618 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4619 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4620 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4621 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4622 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4623 \$1795 \$1773 \$1794 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4624 \$920 \$1773 \$1795 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4625 \$1797 \$1773 \$1796 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4626 \$1798 \$1773 \$1797 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4627 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4628 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4629 \$1799 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4630 \$1800 \$1773 \$1799 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4631 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4632 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4633 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4634 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4635 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4636 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4637 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4638 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4639 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4640 \$1957 \$1730 \$1801 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4641 \$1958 \$1730 \$1957 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4642 \$1802 \$1730 \$1801 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4643 \$1731 \$1730 \$1802 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4644 \$1803 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4645 \$1804 \$1730 \$1803 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4646 \$1960 \$1730 \$1959 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4647 \$1804 \$1730 \$1960 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4648 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4649 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4650 \$1962 \$1730 \$1961 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4651 \$1806 \$1730 \$1962 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4652 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4653 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4654 \$1805 \$1730 \$1731 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4655 \$1806 \$1730 \$1805 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4656 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4657 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4658 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4659 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4660 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4661 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4662 \$1808 \$1730 \$1807 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4663 \$1732 \$1730 \$1808 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4664 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4665 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4666 \$1963 \$1730 \$1807 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4667 \$1964 \$1730 \$1963 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4668 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4669 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4670 \$1809 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4671 \$1810 \$1730 \$1809 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4672 \$1966 \$1730 \$1965 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4673 \$1810 \$1730 \$1966 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4674 \$1811 \$1730 \$1732 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4675 \$1812 \$1730 \$1811 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4676 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4677 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4678 \$1968 \$1730 \$1967 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4679 \$1812 \$1730 \$1968 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4680 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4681 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4682 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4683 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4684 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4685 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4686 \$1969 \$1730 \$1813 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4687 \$1970 \$1730 \$1969 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4688 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4689 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4690 \$1814 \$1730 \$1813 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4691 \$1733 \$1730 \$1814 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4692 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4693 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4694 \$1815 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4695 \$1816 \$1730 \$1815 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4696 \$1972 \$1730 \$1971 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4697 \$1816 \$1730 \$1972 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4698 \$1974 \$1730 \$1973 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4699 \$1818 \$1730 \$1974 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4700 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$4701 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4702 \$1817 \$1730 \$1733 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4703 \$1818 \$1730 \$1817 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4704 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4705 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4706 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4707 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4708 \$1939 \$1773 \$1780 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4709 \$1940 \$1773 \$1939 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4710 \$1942 \$1773 \$1941 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4711 \$1784 \$1773 \$1942 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4712 \$1944 \$1773 \$1943 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4713 \$1786 \$1773 \$1944 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4714 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4715 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4716 \$1945 \$1773 \$1787 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4717 \$1946 \$1773 \$1945 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4718 \$1948 \$1773 \$1947 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4719 \$1791 \$1773 \$1948 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4720 \$1950 \$1773 \$1949 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4721 \$1793 \$1773 \$1950 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4722 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4723 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4724 \$1951 \$1773 \$1794 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4725 \$1952 \$1773 \$1951 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4726 \$1954 \$1773 \$1953 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4727 \$1798 \$1773 \$1954 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4728 \$1956 \$1773 \$1955 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4729 \$1800 \$1773 \$1956 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4730 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4731 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4732 \$2129 \$1773 \$2128 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4733 \$1940 \$1773 \$2129 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4734 \$2130 \$1773 \$1941 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4735 \$2131 \$1773 \$2130 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4736 \$2132 \$1773 \$1943 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4737 \$2133 \$1773 \$2132 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4738 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4739 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4740 \$2135 \$1773 \$2134 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4741 \$1946 \$1773 \$2135 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4742 \$2136 \$1773 \$1947 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4743 \$2137 \$1773 \$2136 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4744 \$2138 \$1773 \$1949 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4745 \$2139 \$1773 \$2138 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4746 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4747 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4748 \$2141 \$1773 \$2140 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4749 \$1952 \$1773 \$2141 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4750 \$2142 \$1773 \$1953 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4751 \$2143 \$1773 \$2142 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4752 \$2144 \$1773 \$1955 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4753 \$2145 \$1773 \$2144 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4754 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4755 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4756 \$2102 \$1730 \$2101 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4757 \$1958 \$1730 \$2102 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4758 \$2103 \$1730 \$1959 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4759 \$2047 \$1730 \$2103 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4760 \$2104 \$1730 \$1961 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4761 \$2105 \$1730 \$2104 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4762 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4763 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4764 \$2107 \$1730 \$2106 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4765 \$1964 \$1730 \$2107 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4766 \$2108 \$1730 \$1965 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4767 \$2048 \$1730 \$2108 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4768 \$2109 \$1730 \$1967 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4769 \$2110 \$1730 \$2109 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4770 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4771 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4772 \$2112 \$1730 \$2111 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4773 \$1970 \$1730 \$2112 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4774 \$2113 \$1730 \$1971 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4775 \$2049 \$1730 \$2113 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4776 \$2114 \$1730 \$1973 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4777 \$2115 \$1730 \$2114 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4778 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4779 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4780 \$2265 \$1773 \$2128 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4781 \$2266 \$1773 \$2265 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4782 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4783 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4784 \$2268 \$1773 \$2267 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4785 \$2133 \$1773 \$2268 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4786 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4787 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4788 \$2269 \$1773 \$2134 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4789 \$2270 \$1773 \$2269 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4790 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4791 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4792 \$2272 \$1773 \$2271 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4793 \$2139 \$1773 \$2272 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4794 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4795 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4796 \$2273 \$1773 \$2140 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4797 \$2274 \$1773 \$2273 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4798 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4799 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4800 \$2276 \$1773 \$2275 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4801 \$2145 \$1773 \$2276 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4802 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4803 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4804 \$2277 \$1730 \$2101 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4805 \$2278 \$1730 \$2277 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4806 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4807 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4808 \$2280 \$1730 \$2279 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4809 \$2105 \$1730 \$2280 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4810 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4811 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4812 \$2281 \$1730 \$2106 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4813 \$2282 \$1730 \$2281 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4814 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4815 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4816 \$2284 \$1730 \$2283 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4817 \$2110 \$1730 \$2284 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4818 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4819 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4820 \$2285 \$1730 \$2111 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4821 \$2286 \$1730 \$2285 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4822 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4823 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4824 \$2288 \$1730 \$2287 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4825 \$2115 \$1730 \$2288 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4826 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4827 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4828 \$2406 \$1773 \$866 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4829 \$1782 \$1773 \$2406 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4830 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4831 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4832 \$2407 \$1773 \$2131 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4833 \$2408 \$1773 \$2407 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4834 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4835 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4836 \$2409 \$1773 \$867 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4837 \$1789 \$1773 \$2409 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4838 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4839 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4840 \$2410 \$1773 \$2137 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4841 \$2411 \$1773 \$2410 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4842 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4843 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4844 \$2412 \$1773 \$868 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4845 \$1796 \$1773 \$2412 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4846 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4847 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4848 \$2413 \$1773 \$2143 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4849 \$2414 \$1773 \$2413 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4850 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4851 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4852 \$2415 \$1730 \$5051 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4853 \$2416 \$1730 \$2415 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4854 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4855 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4856 \$2417 \$1730 \$2442 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4857 \$2047 \$1730 \$2417 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4858 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4859 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4860 \$2418 \$1730 \$5052 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4861 \$2419 \$1730 \$2418 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4862 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4863 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4864 \$2420 \$1730 \$2443 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4865 \$2048 \$1730 \$2420 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4866 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4867 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4868 \$2421 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4869 \$2422 \$1730 \$2421 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4870 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4871 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4872 \$2423 \$1730 \$2444 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4873 \$2049 \$1730 \$2423 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4874 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4875 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4876 \$2608 \$1773 \$2607 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4877 \$2266 \$1773 \$2608 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4878 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4879 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4880 \$2609 \$1773 \$2267 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4881 \$2610 \$1773 \$2609 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4882 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4883 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4884 \$2612 \$1773 \$2611 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4885 \$2270 \$1773 \$2612 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4886 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4887 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4888 \$2613 \$1773 \$2271 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4889 \$2614 \$1773 \$2613 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4890 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4891 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4892 \$2616 \$1773 \$2615 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4893 \$2274 \$1773 \$2616 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4894 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4895 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4896 \$2617 \$1773 \$2275 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4897 \$2618 \$1773 \$2617 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4898 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4899 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4900 \$2584 \$1730 \$2583 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4901 \$2278 \$1730 \$2584 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4902 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4903 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4904 \$2585 \$1730 \$2279 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4905 \$2586 \$1730 \$2585 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4906 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4907 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4908 \$2588 \$1730 \$2587 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4909 \$2282 \$1730 \$2588 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4910 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4911 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4912 \$2589 \$1730 \$2283 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4913 \$2590 \$1730 \$2589 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4914 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4915 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4916 \$2592 \$1730 \$2591 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4917 \$2286 \$1730 \$2592 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4918 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4919 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4920 \$2593 \$1730 \$2287 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4921 \$2594 \$1730 \$2593 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4922 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4923 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4924 \$2745 \$1773 \$2607 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4925 \$2746 \$1773 \$2745 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4926 \$2748 \$1773 \$2747 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4927 \$2408 \$1773 \$2748 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4928 \$2750 \$1773 \$2749 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4929 \$2610 \$1773 \$2750 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4930 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4931 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4932 \$2751 \$1773 \$2611 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4933 \$2752 \$1773 \$2751 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4934 \$2754 \$1773 \$2753 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4935 \$2411 \$1773 \$2754 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4936 \$2756 \$1773 \$2755 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4937 \$2614 \$1773 \$2756 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4938 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4939 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4940 \$2757 \$1773 \$2615 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4941 \$2758 \$1773 \$2757 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4942 \$2760 \$1773 \$2759 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4943 \$2414 \$1773 \$2760 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4944 \$2762 \$1773 \$2761 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4945 \$2618 \$1773 \$2762 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4946 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4947 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4948 \$2763 \$1730 \$2583 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4949 \$2764 \$1730 \$2763 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4950 \$2766 \$1730 \$2765 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4951 \$2442 \$1730 \$2766 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4952 \$2768 \$1730 \$2767 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4953 \$2586 \$1730 \$2768 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4954 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4955 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4956 \$2769 \$1730 \$2587 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4957 \$2770 \$1730 \$2769 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4958 \$2772 \$1730 \$2771 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4959 \$2443 \$1730 \$2772 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4960 \$2774 \$1730 \$2773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4961 \$2590 \$1730 \$2774 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4962 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4963 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4964 \$2775 \$1730 \$2591 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4965 \$2776 \$1730 \$2775 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4966 \$2778 \$1730 \$2777 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4967 \$2444 \$1730 \$2778 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4968 \$2780 \$1730 \$2779 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4969 \$2594 \$1730 \$2780 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4970 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4971 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4972 \$2900 \$1773 \$2899 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4973 \$2746 \$1773 \$2900 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4974 \$2901 \$1773 \$2747 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4975 \$2902 \$1773 \$2901 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4976 \$2903 \$1773 \$2749 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4977 \$2904 \$1773 \$2903 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4978 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4979 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4980 \$2906 \$1773 \$2905 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4981 \$2752 \$1773 \$2906 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4982 \$2907 \$1773 \$2753 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4983 \$2908 \$1773 \$2907 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4984 \$2909 \$1773 \$2755 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4985 \$2910 \$1773 \$2909 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4986 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4987 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4988 \$2912 \$1773 \$2911 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4989 \$2758 \$1773 \$2912 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4990 \$2913 \$1773 \$2759 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4991 \$2914 \$1773 \$2913 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4992 \$2915 \$1773 \$2761 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4993 \$2916 \$1773 \$2915 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4994 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4995 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4996 \$2918 \$1730 \$2917 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4997 \$2764 \$1730 \$2918 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$4998 \$2919 \$1730 \$2765 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$4999 \$2920 \$1730 \$2919 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5000 \$2921 \$1730 \$2767 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5001 \$2922 \$1730 \$2921 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5002 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5003 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5004 \$2924 \$1730 \$2923 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5005 \$2770 \$1730 \$2924 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5006 \$2925 \$1730 \$2771 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5007 \$2926 \$1730 \$2925 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5008 \$2927 \$1730 \$2773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5009 \$2928 \$1730 \$2927 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5010 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5011 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5012 \$2930 \$1730 \$2929 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5013 \$2776 \$1730 \$2930 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5014 \$2931 \$1730 \$2777 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5015 \$2932 \$1730 \$2931 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5016 \$2933 \$1730 \$2779 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5017 \$2934 \$1730 \$2933 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5018 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5019 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5020 \$3052 \$1773 \$2899 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5021 \$3053 \$1773 \$3052 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5022 \$3054 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5023 \$2902 \$1773 \$3054 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5024 \$3055 \$1773 \$3053 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5025 \$2904 \$1773 \$3055 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5026 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5027 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5028 \$3056 \$1773 \$2905 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5029 \$3057 \$1773 \$3056 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5030 \$3058 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5031 \$2908 \$1773 \$3058 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5032 \$3059 \$1773 \$3057 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5033 \$2910 \$1773 \$3059 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5034 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5035 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5036 \$3060 \$1773 \$2911 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5037 \$3061 \$1773 \$3060 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5038 \$3062 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5039 \$2914 \$1773 \$3062 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5040 \$3063 \$1773 \$3061 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5041 \$2916 \$1773 \$3063 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5042 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5043 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5044 \$3064 \$1730 \$2917 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5045 \$3065 \$1730 \$3064 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5046 \$3066 \$1730 \$2416 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5047 \$2920 \$1730 \$3066 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5048 \$3067 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5049 \$2922 \$1730 \$3067 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5050 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5051 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5052 \$3068 \$1730 \$2923 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5053 \$3069 \$1730 \$3068 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5054 \$3070 \$1730 \$2419 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5055 \$2926 \$1730 \$3070 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5056 \$3071 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5057 \$2928 \$1730 \$3071 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5058 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5059 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5060 \$3072 \$1730 \$2929 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5061 CMOUTN \$1730 \$3072 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5062 \$3074 \$1730 \$2422 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5063 \$2932 \$1730 \$3074 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5064 \$3075 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5065 \$2934 \$1730 \$3075 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5066 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5067 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5068 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5069 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5070 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5071 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5072 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5073 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5074 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5075 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5076 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5077 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5078 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5079 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5080 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5081 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5082 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5083 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5084 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5085 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5086 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5087 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5088 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5089 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5090 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5091 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5092 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5093 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5094 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5095 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5096 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5097 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5098 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5099 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5100 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5101 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5102 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5103 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5104 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5105 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5106 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5107 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5108 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5109 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5110 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5111 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5112 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5113 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5114 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5115 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5116 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5117 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5118 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5119 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5120 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5121 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5122 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5123 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5124 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5125 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5126 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5127 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5128 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5129 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5130 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5131 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5132 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5133 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5134 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5135 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5136 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5137 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5138 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5139 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5140 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5141 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5142 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5143 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5144 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5145 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5146 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5147 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5148 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5149 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5150 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5151 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5152 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5153 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5154 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5155 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5156 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5157 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5158 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5159 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5160 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5161 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5162 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5163 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5164 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5165 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5166 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5167 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5168 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5169 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5170 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5171 \$3166 ISBCS ISBCS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5172 VSS ISBCS \$3166 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5173 \$3252 ISBCS \$1573 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5174 VSS ISBCS \$3252 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5175 \$3167 ISBCS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5176 \$1574 ISBCS \$3167 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5177 \$3253 ISBCS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5178 \$4093 ISBCS \$3253 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5179 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5180 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5181 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5182 \$3398 \$1773 \$3397 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5183 \$922 \$1773 \$3398 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5184 \$3400 \$1773 \$3399 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5185 \$3401 \$1773 \$3400 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5186 \$3402 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5187 \$3403 \$1773 \$3402 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5188 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5189 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5190 \$3405 \$1773 \$3404 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5191 \$924 \$1773 \$3405 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5192 \$3407 \$1773 \$3406 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5193 \$3408 \$1773 \$3407 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5194 \$3409 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5195 \$3410 \$1773 \$3409 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5196 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5197 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5198 \$3412 \$1773 \$3411 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5199 VSS \$1773 \$3412 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5200 \$3414 \$1773 \$3413 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5201 \$3415 \$1773 \$3414 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5202 \$3416 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5203 \$3417 \$1773 \$3416 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5204 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5205 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5206 \$3419 \$1730 \$3418 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5207 \$3376 \$1730 \$3419 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5208 \$3420 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5209 \$3421 \$1730 \$3420 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5210 \$3422 \$1730 \$3376 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5211 \$3423 \$1730 \$3422 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5212 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5213 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5214 \$3425 \$1730 \$3424 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5215 \$3377 \$1730 \$3425 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5216 \$3426 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5217 \$3427 \$1730 \$3426 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5218 \$3428 \$1730 \$3377 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5219 \$3429 \$1730 \$3428 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5220 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5221 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5222 \$3431 \$1730 \$3430 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5223 \$3378 \$1730 \$3431 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5224 \$3432 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5225 \$3433 \$1730 \$3432 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5226 \$3434 \$1730 \$3378 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5227 \$3435 \$1730 \$3434 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5228 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5229 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5230 \$3332 ISBCS \$1573 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5231 VSS ISBCS \$3332 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5232 \$3333 ISBCS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5233 \$4093 ISBCS \$3333 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5234 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5235 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5236 \$3569 \$1773 \$3397 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5237 \$3570 \$1773 \$3569 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5238 \$3572 \$1773 \$3571 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5239 \$3401 \$1773 \$3572 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5240 \$3574 \$1773 \$3573 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5241 \$3403 \$1773 \$3574 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5242 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5243 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5244 \$3575 \$1773 \$3404 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5245 \$3576 \$1773 \$3575 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5246 \$3578 \$1773 \$3577 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5247 \$3408 \$1773 \$3578 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5248 \$3580 \$1773 \$3579 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5249 \$3410 \$1773 \$3580 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5250 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5251 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5252 \$3581 \$1773 \$3411 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5253 \$3582 \$1773 \$3581 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5254 \$3584 \$1773 \$3583 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5255 \$3415 \$1773 \$3584 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5256 \$3586 \$1773 \$3585 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5257 \$3417 \$1773 \$3586 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5258 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5259 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5260 \$3587 \$1730 \$3418 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5261 \$3588 \$1730 \$3587 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5262 \$3590 \$1730 \$3589 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5263 \$3421 \$1730 \$3590 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5264 \$3592 \$1730 \$3591 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5265 \$3423 \$1730 \$3592 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5266 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5267 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5268 \$3593 \$1730 \$3424 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5269 \$3594 \$1730 \$3593 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5270 \$3596 \$1730 \$3595 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5271 \$3427 \$1730 \$3596 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5272 \$3598 \$1730 \$3597 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5273 \$3429 \$1730 \$3598 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5274 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5275 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5276 \$3599 \$1730 \$3430 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5277 \$3600 \$1730 \$3599 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5278 \$3602 \$1730 \$3601 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5279 \$3433 \$1730 \$3602 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5280 \$3604 \$1730 \$3603 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5281 \$3435 \$1730 \$3604 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5282 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5283 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5284 \$3477 ISBCS \$1574 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5285 VSS ISBCS \$3477 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5286 \$3478 ISBCS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5287 ISBCS ISBCS \$3478 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5288 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5289 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5290 \$3729 \$1773 \$3728 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5291 \$3570 \$1773 \$3729 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5292 \$3730 \$1773 \$3571 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5293 \$3731 \$1773 \$3730 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5294 \$3732 \$1773 \$3573 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5295 \$3733 \$1773 \$3732 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5296 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5297 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5298 \$3735 \$1773 \$3734 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5299 \$3576 \$1773 \$3735 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5300 \$3736 \$1773 \$3577 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5301 \$3737 \$1773 \$3736 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5302 \$3738 \$1773 \$3579 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5303 \$3739 \$1773 \$3738 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5304 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5305 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5306 \$3741 \$1773 \$3740 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5307 \$3582 \$1773 \$3741 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5308 \$3742 \$1773 \$3583 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5309 \$3743 \$1773 \$3742 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5310 \$3744 \$1773 \$3585 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5311 \$3745 \$1773 \$3744 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5312 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5313 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5314 \$3747 \$1730 \$3746 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5315 \$3588 \$1730 \$3747 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5316 \$3748 \$1730 \$3589 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5317 \$3642 \$1730 \$3748 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5318 \$3749 \$1730 \$3591 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5319 \$3750 \$1730 \$3749 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5320 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5321 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5322 \$3752 \$1730 \$3751 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5323 \$3594 \$1730 \$3752 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5324 \$3753 \$1730 \$3595 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5325 \$3643 \$1730 \$3753 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5326 \$3754 \$1730 \$3597 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5327 \$3755 \$1730 \$3754 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5328 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5329 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5330 \$3757 \$1730 \$3756 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5331 \$3600 \$1730 \$3757 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5332 \$3758 \$1730 \$3601 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5333 \$3644 \$1730 \$3758 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5334 \$3759 \$1730 \$3603 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5335 \$3760 \$1730 \$3759 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5336 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5337 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5338 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5339 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5340 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5341 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5342 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5343 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5344 \$3901 \$1773 \$3728 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5345 \$3902 \$1773 \$3901 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5346 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5347 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5348 \$3904 \$1773 \$3903 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5349 \$3733 \$1773 \$3904 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5350 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5351 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5352 \$3905 \$1773 \$3734 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5353 \$3906 \$1773 \$3905 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5354 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5355 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5356 \$3908 \$1773 \$3907 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5357 \$3739 \$1773 \$3908 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5358 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5359 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5360 \$3909 \$1773 \$3740 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5361 \$3910 \$1773 \$3909 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5362 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5363 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5364 \$3912 \$1773 \$3911 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5365 \$3745 \$1773 \$3912 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5366 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5367 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5368 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5369 \$4074 \$1730 \$5048 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5370 \$4075 \$1730 \$4074 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5371 \$3913 \$1730 \$3746 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5372 \$3914 \$1730 \$3913 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5373 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5374 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5375 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5376 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5377 \$4077 \$1730 \$4076 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5378 \$3642 \$1730 \$4077 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5379 \$3916 \$1730 \$3915 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5380 \$3750 \$1730 \$3916 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5381 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5382 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5383 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5384 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5385 \$4078 \$1730 \$5049 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5386 \$4079 \$1730 \$4078 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5387 \$3917 \$1730 \$3751 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5388 \$3918 \$1730 \$3917 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5389 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5390 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5391 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5392 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5393 \$3920 \$1730 \$3919 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5394 \$3755 \$1730 \$3920 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5395 \$4081 \$1730 \$4080 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5396 \$3643 \$1730 \$4081 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5397 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5398 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5399 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5400 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5401 \$4082 \$1730 \$5050 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5402 \$4083 \$1730 \$4082 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5403 \$3921 \$1730 \$3756 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5404 \$3922 \$1730 \$3921 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5405 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5406 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5407 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5408 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5409 \$4085 \$1730 \$4084 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5410 \$3644 \$1730 \$4085 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5411 \$3924 \$1730 \$3923 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5412 \$3760 \$1730 \$3924 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5413 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5414 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5415 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5416 \$4065 \$1773 \$869 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5417 \$3399 \$1773 \$4065 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5418 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5419 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5420 \$4066 \$1773 \$3731 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5421 \$4067 \$1773 \$4066 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5422 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5423 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5424 \$4068 \$1773 \$870 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5425 \$3406 \$1773 \$4068 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5426 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5427 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5428 \$4069 \$1773 \$3737 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5429 \$4070 \$1773 \$4069 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5430 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5431 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5432 \$4071 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5433 \$3413 \$1773 \$4071 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5434 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5435 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5436 \$4072 \$1773 \$3743 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5437 \$4073 \$1773 \$4072 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5438 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5439 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5440 \$4225 \$1773 \$4224 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5441 \$3902 \$1773 \$4225 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5442 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5443 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5444 \$4226 \$1773 \$3903 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5445 \$4227 \$1773 \$4226 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5446 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5447 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5448 \$4229 \$1773 \$4228 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5449 \$3906 \$1773 \$4229 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5450 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5451 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5452 \$4230 \$1773 \$3907 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5453 \$4231 \$1773 \$4230 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5454 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5455 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5456 \$4233 \$1773 \$4232 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5457 \$3910 \$1773 \$4233 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5458 VSS \$1773 \$1773 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5459 \$1773 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5460 \$4234 \$1773 \$3911 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5461 \$4235 \$1773 \$4234 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5462 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5463 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5464 \$4237 \$1730 \$4236 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5465 \$3914 \$1730 \$4237 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5466 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5467 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5468 \$4238 \$1730 \$3915 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5469 \$4239 \$1730 \$4238 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5470 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5471 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5472 \$4241 \$1730 \$4240 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5473 \$3918 \$1730 \$4241 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5474 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5475 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5476 \$4242 \$1730 \$3919 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5477 \$4243 \$1730 \$4242 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5478 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5479 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5480 \$4245 \$1730 \$4244 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5481 \$3922 \$1730 \$4245 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5482 VSS \$1730 \$1730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5483 \$1730 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5484 \$4246 \$1730 \$3923 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5485 \$4247 \$1730 \$4246 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5486 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5487 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5488 \$4407 \$1773 \$4224 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5489 \$4408 \$1773 \$4407 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5490 \$4410 \$1773 \$4409 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5491 \$4067 \$1773 \$4410 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5492 \$4412 \$1773 \$4411 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5493 \$4227 \$1773 \$4412 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5494 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5495 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5496 \$4413 \$1773 \$4228 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5497 \$4414 \$1773 \$4413 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5498 \$4416 \$1773 \$4415 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5499 \$4070 \$1773 \$4416 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5500 \$4418 \$1773 \$4417 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5501 \$4231 \$1773 \$4418 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5502 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5503 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5504 \$4419 \$1773 \$4232 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5505 \$4420 \$1773 \$4419 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5506 \$4422 \$1773 \$4421 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5507 \$4073 \$1773 \$4422 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5508 \$4424 \$1773 \$4423 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5509 \$4235 \$1773 \$4424 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5510 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5511 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5512 \$4425 \$1730 \$4236 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5513 \$4426 \$1730 \$4425 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5514 \$4428 \$1730 \$4427 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5515 \$4076 \$1730 \$4428 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5516 \$4430 \$1730 \$4429 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5517 \$4239 \$1730 \$4430 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5518 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5519 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5520 \$4431 \$1730 \$4240 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5521 \$4432 \$1730 \$4431 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5522 \$4434 \$1730 \$4433 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5523 \$4080 \$1730 \$4434 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5524 \$4436 \$1730 \$4435 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5525 \$4243 \$1730 \$4436 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5526 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5527 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5528 \$4437 \$1730 \$4244 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5529 \$4438 \$1730 \$4437 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5530 \$4440 \$1730 \$4439 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5531 \$4084 \$1730 \$4440 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5532 \$4442 \$1730 \$4441 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5533 \$4247 \$1730 \$4442 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5534 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5535 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5536 \$4573 \$1773 \$4572 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5537 \$4408 \$1773 \$4573 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5538 \$4574 \$1773 \$4409 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5539 \$4575 \$1773 \$4574 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5540 \$4576 \$1773 \$4411 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5541 \$4577 \$1773 \$4576 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5542 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5543 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5544 \$4579 \$1773 \$4578 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5545 \$4414 \$1773 \$4579 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5546 \$4580 \$1773 \$4415 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5547 \$4581 \$1773 \$4580 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5548 \$4582 \$1773 \$4417 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5549 \$4583 \$1773 \$4582 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5550 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5551 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5552 \$4585 \$1773 \$4584 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5553 \$4420 \$1773 \$4585 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5554 \$4586 \$1773 \$4421 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5555 \$4587 \$1773 \$4586 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5556 \$4588 \$1773 \$4423 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5557 \$4589 \$1773 \$4588 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5558 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5559 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5560 \$4591 \$1730 \$4590 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5561 \$4426 \$1730 \$4591 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5562 \$4592 \$1730 \$4427 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5563 \$4593 \$1730 \$4592 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5564 \$4594 \$1730 \$4429 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5565 \$4595 \$1730 \$4594 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5566 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5567 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5568 \$4597 \$1730 \$4596 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5569 \$4432 \$1730 \$4597 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5570 \$4598 \$1730 \$4433 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5571 \$4599 \$1730 \$4598 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5572 \$4600 \$1730 \$4435 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5573 \$4601 \$1730 \$4600 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5574 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5575 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5576 \$4603 \$1730 \$4602 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5577 \$4438 \$1730 \$4603 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5578 \$4604 \$1730 \$4439 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5579 \$4605 \$1730 \$4604 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5580 \$4606 \$1730 \$4441 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5581 \$4607 \$1730 \$4606 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5582 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5583 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5584 \$4713 \$1773 \$4572 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5585 \$4714 \$1773 \$4713 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5586 \$4715 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5587 \$4575 \$1773 \$4715 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5588 \$4716 \$1773 \$4714 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5589 \$4577 \$1773 \$4716 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5590 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5591 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5592 \$4717 \$1773 \$4578 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5593 \$4718 \$1773 \$4717 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5594 \$4719 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5595 \$4581 \$1773 \$4719 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5596 \$4720 \$1773 \$4718 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5597 \$4583 \$1773 \$4720 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5598 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5599 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5600 \$4721 \$1773 \$4584 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5601 \$4722 \$1773 \$4721 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5602 \$4723 \$1773 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5603 \$4587 \$1773 \$4723 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5604 \$4724 \$1773 \$4722 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5605 \$4589 \$1773 \$4724 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5606 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5607 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5608 \$4725 \$1730 \$4590 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5609 \$4726 \$1730 \$4725 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5610 \$4727 \$1730 \$4075 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5611 \$4593 \$1730 \$4727 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5612 \$4728 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5613 \$4595 \$1730 \$4728 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5614 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5615 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5616 \$4729 \$1730 \$4596 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5617 \$4730 \$1730 \$4729 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5618 \$4731 \$1730 \$4079 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5619 \$4599 \$1730 \$4731 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5620 \$4732 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5621 \$4601 \$1730 \$4732 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5622 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5623 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5624 \$4733 \$1730 \$4602 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5625 \$4734 \$1730 \$4733 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5626 \$4735 \$1730 \$4083 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5627 \$4605 \$1730 \$4735 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5628 \$4736 \$1730 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5629 \$4607 \$1730 \$4736 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5630 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5631 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5632 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5633 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5634 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5635 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5636 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5637 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5638 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5639 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5640 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5641 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5642 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5643 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5644 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5645 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5646 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5647 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5648 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5649 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5650 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5651 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5652 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5653 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5654 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5655 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5656 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5657 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5658 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5659 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5660 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5661 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5662 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5663 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5664 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5665 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5666 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5667 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5668 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5669 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5670 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5671 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5672 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5673 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5674 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5675 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5676 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5677 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5678 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5679 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5680 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5681 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5682 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5683 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5684 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5685 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5686 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5687 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5688 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5689 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5690 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5691 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5692 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5693 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5694 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5695 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5696 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5697 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5698 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5699 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5700 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5701 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5702 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5703 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5704 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5705 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5706 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5707 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5708 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5709 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5710 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5711 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5712 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5713 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5714 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5715 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5716 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5717 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5718 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5719 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5720 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5721 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5722 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5723 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5724 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5725 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5726 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5727 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5728 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5729 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5730 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5731 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5732 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5733 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5734 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5735 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5736 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5737 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5738 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5739 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5740 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5741 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5742 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5743 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5744 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5745 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5746 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5747 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5748 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5749 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5750 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5751 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5752 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5753 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5754 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5755 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5756 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5757 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5758 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5759 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5760 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5761 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5762 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5763 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5764 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5765 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5766 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5767 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5768 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5769 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5770 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5771 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5772 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5773 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5774 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5775 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5776 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5777 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5778 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5779 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5780 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5781 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5782 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5783 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5784 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5785 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5786 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5787 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5788 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5789 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5790 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5791 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5792 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5793 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5794 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5795 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5796 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5797 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5798 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5799 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5800 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5801 \$5074 \$5113 \$5073 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5802 \$5048 \$5113 \$5074 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5803 \$5075 \$4726 \$5048 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5804 \$4973 \$4726 \$5075 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5805 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5806 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5807 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5808 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5809 \$5077 \$4973 \$5076 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5810 \$5113 \$4973 \$5077 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5811 \$5078 \$4973 \$5113 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5812 \$5183 \$4973 \$5078 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5813 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5814 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5815 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5816 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5817 \$5079 \$5114 \$5114 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5818 VSS \$5114 \$5079 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5819 \$5080 \$5114 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5820 \$5850 \$5114 \$5080 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5821 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5822 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5823 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5824 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5825 \$5082 \$5115 \$5081 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5826 \$5049 \$5115 \$5082 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5827 \$5083 \$4730 \$5049 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5828 \$4974 \$4730 \$5083 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5829 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5830 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5831 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5832 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5833 \$5085 \$4974 \$5084 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5834 \$5115 \$4974 \$5085 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5835 \$5086 \$4974 \$5115 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5836 \$5184 \$4974 \$5086 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5837 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5838 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5839 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5840 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5841 \$5087 \$5116 \$5116 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5842 VSS \$5116 \$5087 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5843 \$5088 \$5116 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5844 \$5851 \$5116 \$5088 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5845 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5846 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5847 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5848 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5849 \$5090 \$5117 \$5089 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5850 \$5050 \$5117 \$5090 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5851 \$5091 \$4734 \$5050 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5852 \$4975 \$4734 \$5091 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5853 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5854 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5855 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5856 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5857 \$5093 \$4975 \$5092 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5858 \$5117 \$4975 \$5093 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5859 \$5094 \$4975 \$5117 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5860 \$5185 \$4975 \$5094 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5861 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5862 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5863 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5864 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5865 \$5095 \$5118 \$5118 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5866 VSS \$5118 \$5095 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5867 \$5096 \$5118 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5868 \$5852 \$5118 \$5096 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5869 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5870 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5871 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5872 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5873 \$5098 \$5119 \$5097 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5874 \$5051 \$5119 \$5098 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5875 \$5099 \$3065 \$5051 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5876 \$4976 \$3065 \$5099 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5877 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5878 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5879 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5880 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5881 \$5101 \$4976 \$5100 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5882 \$5119 \$4976 \$5101 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5883 \$5102 \$4976 \$5119 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5884 \$5186 \$4976 \$5102 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5885 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5886 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5887 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5888 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5889 \$5103 \$5120 \$5120 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5890 VSS \$5120 \$5103 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5891 \$5104 \$5120 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5892 \$5853 \$5120 \$5104 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5893 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5894 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5895 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5896 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5897 \$5106 \$5121 \$5105 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5898 \$5052 \$5121 \$5106 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5899 \$5107 \$3069 \$5052 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5900 \$4977 \$3069 \$5107 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5901 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5902 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5903 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5904 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5905 \$5109 \$4977 \$5108 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5906 \$5121 \$4977 \$5109 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5907 \$5110 \$4977 \$5121 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5908 \$5187 \$4977 \$5110 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5909 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5910 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5911 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5912 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5913 \$5111 \$5122 \$5122 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5914 VSS \$5122 \$5111 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5915 \$5112 \$5122 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5916 \$5854 \$5122 \$5112 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5917 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5918 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5919 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5920 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5921 \$5258 \$4726 \$4973 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5922 \$5048 \$4726 \$5258 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5923 \$5259 \$5113 \$5048 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5924 \$5073 \$5113 \$5259 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5925 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5926 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5927 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5928 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5929 \$5260 \$4973 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5930 \$4726 \$4973 \$5260 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5931 \$5261 \$4973 \$4726 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5932 VDD \$4973 \$5261 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5933 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5934 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5935 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5936 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5937 \$5262 \$5114 \$5850 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5938 VSS \$5114 \$5262 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5939 \$5263 \$5114 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5940 \$5114 \$5114 \$5263 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5941 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5942 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5943 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5944 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5945 \$5264 \$4730 \$4974 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5946 \$5049 \$4730 \$5264 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5947 \$5265 \$5115 \$5049 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5948 \$5081 \$5115 \$5265 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5949 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5950 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5951 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5952 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5953 \$5266 \$4974 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5954 \$4730 \$4974 \$5266 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5955 \$5267 \$4974 \$4730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5956 VDD \$4974 \$5267 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5957 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5958 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5959 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5960 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5961 \$5268 \$5116 \$5851 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5962 VSS \$5116 \$5268 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5963 \$5269 \$5116 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5964 \$5116 \$5116 \$5269 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5965 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5966 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5967 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5968 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5969 \$5270 \$4734 \$4975 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5970 \$5050 \$4734 \$5270 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5971 \$5271 \$5117 \$5050 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5972 \$5089 \$5117 \$5271 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5973 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5974 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5975 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5976 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5977 \$5272 \$4975 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5978 \$4734 \$4975 \$5272 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5979 \$5273 \$4975 \$4734 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5980 VDD \$4975 \$5273 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5981 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5982 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5983 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5984 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5985 \$5274 \$5118 \$5852 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5986 VSS \$5118 \$5274 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5987 \$5275 \$5118 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5988 \$5118 \$5118 \$5275 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5989 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5990 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5991 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5992 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5993 \$5276 \$3065 \$4976 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5994 \$5051 \$3065 \$5276 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5995 \$5277 \$5119 \$5051 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$5996 \$5097 \$5119 \$5277 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$5997 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5998 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$5999 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6000 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6001 \$5278 \$4976 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6002 \$3065 \$4976 \$5278 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6003 \$5279 \$4976 \$3065 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6004 VDD \$4976 \$5279 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6005 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6006 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6007 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6008 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6009 \$5280 \$5120 \$5853 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6010 VSS \$5120 \$5280 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6011 \$5281 \$5120 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6012 \$5120 \$5120 \$5281 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6013 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6014 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6015 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6016 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6017 \$5282 \$3069 \$4977 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6018 \$5052 \$3069 \$5282 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6019 \$5283 \$5121 \$5052 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6020 \$5105 \$5121 \$5283 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6021 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6022 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6023 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6024 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6025 \$5284 \$4977 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6026 \$3069 \$4977 \$5284 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6027 \$5285 \$4977 \$3069 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6028 VDD \$4977 \$5285 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6029 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6030 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6031 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6032 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6033 \$5286 \$5122 \$5854 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6034 VSS \$5122 \$5286 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6035 \$5287 \$5122 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6036 \$5122 \$5122 \$5287 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6037 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6038 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6039 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6040 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6041 \$5378 \$5113 \$5073 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6042 \$5048 \$5113 \$5378 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6043 \$5379 \$4726 \$5048 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6044 \$4973 \$4726 \$5379 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6045 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6046 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6047 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6048 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6049 \$5380 \$4973 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6050 \$4726 \$4973 \$5380 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6051 \$5381 \$4973 \$4726 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6052 VDD \$4973 \$5381 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6053 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6054 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6055 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6056 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6057 \$5382 \$5114 \$5114 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6058 VSS \$5114 \$5382 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6059 \$5383 \$5114 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6060 \$5850 \$5114 \$5383 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6061 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6062 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6063 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6064 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6065 \$5384 \$5115 \$5081 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6066 \$5049 \$5115 \$5384 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6067 \$5385 \$4730 \$5049 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6068 \$4974 \$4730 \$5385 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6069 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6070 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6071 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6072 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6073 \$5386 \$4974 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6074 \$4730 \$4974 \$5386 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6075 \$5387 \$4974 \$4730 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6076 VDD \$4974 \$5387 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6077 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6078 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6079 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6080 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6081 \$5388 \$5116 \$5116 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6082 VSS \$5116 \$5388 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6083 \$5389 \$5116 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6084 \$5851 \$5116 \$5389 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6085 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6086 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6087 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6088 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6089 \$5390 \$5117 \$5089 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6090 \$5050 \$5117 \$5390 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6091 \$5391 \$4734 \$5050 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6092 \$4975 \$4734 \$5391 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6093 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6094 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6095 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6096 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6097 \$5392 \$4975 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6098 \$4734 \$4975 \$5392 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6099 \$5393 \$4975 \$4734 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6100 VDD \$4975 \$5393 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6101 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6102 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6103 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6104 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6105 \$5394 \$5118 \$5118 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6106 VSS \$5118 \$5394 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6107 \$5395 \$5118 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6108 \$5852 \$5118 \$5395 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6109 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6110 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6111 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6112 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6113 \$5396 \$5119 \$5097 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6114 \$5051 \$5119 \$5396 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6115 \$5397 \$3065 \$5051 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6116 \$4976 \$3065 \$5397 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6117 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6118 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6119 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6120 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6121 \$5398 \$4976 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6122 \$3065 \$4976 \$5398 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6123 \$5399 \$4976 \$3065 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6124 VDD \$4976 \$5399 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6125 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6126 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6127 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6128 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6129 \$5400 \$5120 \$5120 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6130 VSS \$5120 \$5400 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6131 \$5401 \$5120 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6132 \$5853 \$5120 \$5401 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6133 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6134 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6135 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6136 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6137 \$5402 \$5121 \$5105 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6138 \$5052 \$5121 \$5402 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6139 \$5403 \$3069 \$5052 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6140 \$4977 \$3069 \$5403 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6141 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6142 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6143 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6144 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6145 \$5404 \$4977 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6146 \$3069 \$4977 \$5404 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6147 \$5405 \$4977 \$3069 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6148 VDD \$4977 \$5405 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6149 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6150 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6151 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6152 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6153 \$5406 \$5122 \$5122 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6154 VSS \$5122 \$5406 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6155 \$5407 \$5122 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6156 \$5854 \$5122 \$5407 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6157 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6158 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6159 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6160 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6161 \$5523 \$4726 \$4973 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6162 \$5048 \$4726 \$5523 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6163 \$5524 \$5113 \$5048 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6164 \$5073 \$5113 \$5524 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6165 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6166 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6167 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6168 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6169 \$5525 \$4973 \$5183 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6170 \$5113 \$4973 \$5525 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6171 \$5526 \$4973 \$5113 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6172 \$5076 \$4973 \$5526 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6173 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6174 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6175 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6176 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6177 \$5527 \$5114 \$5850 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6178 VSS \$5114 \$5527 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6179 \$5528 \$5114 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6180 \$5114 \$5114 \$5528 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6181 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6182 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6183 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6184 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6185 \$5529 \$4730 \$4974 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6186 \$5049 \$4730 \$5529 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6187 \$5530 \$5115 \$5049 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6188 \$5081 \$5115 \$5530 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6189 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6190 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6191 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6192 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6193 \$5531 \$4974 \$5184 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6194 \$5115 \$4974 \$5531 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6195 \$5532 \$4974 \$5115 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6196 \$5084 \$4974 \$5532 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6197 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6198 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6199 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6200 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6201 \$5533 \$5116 \$5851 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6202 VSS \$5116 \$5533 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6203 \$5534 \$5116 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6204 \$5116 \$5116 \$5534 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6205 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6206 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6207 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6208 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6209 \$5535 \$4734 \$4975 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6210 \$5050 \$4734 \$5535 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6211 \$5536 \$5117 \$5050 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6212 \$5089 \$5117 \$5536 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6213 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6214 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6215 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6216 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6217 \$5537 \$4975 \$5185 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6218 \$5117 \$4975 \$5537 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6219 \$5538 \$4975 \$5117 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6220 \$5092 \$4975 \$5538 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6221 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6222 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6223 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6224 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6225 \$5539 \$5118 \$5852 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6226 VSS \$5118 \$5539 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6227 \$5540 \$5118 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6228 \$5118 \$5118 \$5540 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6229 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6230 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6231 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6232 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6233 \$5541 \$3065 \$4976 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6234 \$5051 \$3065 \$5541 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6235 \$5542 \$5119 \$5051 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6236 \$5097 \$5119 \$5542 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6237 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6238 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6239 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6240 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6241 \$5543 \$4976 \$5186 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6242 \$5119 \$4976 \$5543 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6243 \$5544 \$4976 \$5119 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6244 \$5100 \$4976 \$5544 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6245 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6246 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6247 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6248 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6249 \$5545 \$5120 \$5853 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6250 VSS \$5120 \$5545 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6251 \$5546 \$5120 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6252 \$5120 \$5120 \$5546 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6253 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6254 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6255 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6256 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6257 \$5547 \$3069 \$4977 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6258 \$5052 \$3069 \$5547 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6259 \$5548 \$5121 \$5052 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6260 \$5105 \$5121 \$5548 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6261 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6262 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6263 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6264 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6265 \$5549 \$4977 \$5187 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6266 \$5121 \$4977 \$5549 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6267 \$5550 \$4977 \$5121 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6268 \$5108 \$4977 \$5550 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6269 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6270 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6271 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6272 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6273 \$5551 \$5122 \$5854 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6274 VSS \$5122 \$5551 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6275 \$5552 \$5122 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6276 \$5122 \$5122 \$5552 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6277 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6278 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6279 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6280 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6281 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6282 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6283 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6284 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6285 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6286 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6287 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6288 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6289 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6290 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6291 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6292 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6293 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6294 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6295 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6296 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6297 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6298 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6299 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6300 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6301 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6302 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6303 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6304 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6305 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6306 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6307 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6308 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6309 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6310 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6311 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6312 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6313 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6314 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6315 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6316 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6317 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6318 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6319 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6320 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6321 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6322 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6323 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6324 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6325 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6326 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6327 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6328 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6329 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6330 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6331 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6332 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6333 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6334 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6335 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6336 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6337 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6338 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6339 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6340 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6341 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6342 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6343 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6344 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6345 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6346 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6347 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6348 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6349 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6350 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6351 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6352 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6353 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6354 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6355 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6356 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6357 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6358 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6359 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6360 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6361 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6362 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6363 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6364 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6365 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6366 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6367 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6368 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6369 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6370 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6371 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6372 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6373 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6374 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6375 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6376 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6377 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6378 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6379 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6380 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6381 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6382 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6383 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6384 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6385 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6386 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6387 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6388 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6389 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6390 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6391 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6392 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6393 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6394 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6395 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6396 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6397 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6398 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6399 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6400 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6401 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6402 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6403 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6404 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6405 \$9355 ISBCS2 \$8551 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6406 \$9355 ISBCS2 \$10007 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6407 \$7676 ISBCS2 \$8551 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6408 \$7676 ISBCS2 VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6409 ISBCS2 ISBCS2 VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6410 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6411 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6412 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6413 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6414 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6415 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6416 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6417 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6418 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6419 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6420 AVSS \$8587 \$8587 VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P
+ PS=5.72U PD=3.05U
M$6421 \$8587 \$8587 AVSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P
+ PS=3.05U PD=5.72U
M$6422 AVSS \$8587 \$8078 VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P
+ PS=5.72U PD=3.05U
M$6423 \$8078 \$8587 AVSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P
+ PS=3.05U PD=5.72U
M$6424 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$6425 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$6426 AVSS \$8587 \$8078 VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P
+ PS=5.72U PD=3.05U
M$6427 \$8078 \$8587 AVSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P
+ PS=3.05U PD=5.72U
M$6428 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$6429 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$6430 AVSS \$8587 \$8587 VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P
+ PS=5.72U PD=3.05U
M$6431 \$8587 \$8587 AVSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P
+ PS=3.05U PD=5.72U
M$6432 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6433 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6434 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6435 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6436 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6437 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6438 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6439 \$10416 \$9382 \$9382 VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P
+ PS=3.62U PD=2U
M$6440 \$9871 \$9382 \$10416 VSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U
+ PD=3.62U
M$6441 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P PS=3.62U
+ PD=2U
M$6442 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U
+ PD=3.62U
M$6443 \$9870 \$9382 \$9356 VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P
+ PS=3.62U PD=2U
M$6444 \$9871 \$9382 \$9870 VSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U
+ PD=3.62U
M$6445 \$9357 \$9382 \$9356 VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P
+ PS=3.62U PD=2U
M$6446 AVSS \$9382 \$9357 VSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U
+ PD=3.62U
M$6447 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6448 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6449 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6450 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6451 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6452 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6453 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6454 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6455 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6456 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6457 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6458 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6459 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6460 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6461 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6462 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6463 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6464 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6465 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6466 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6467 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6468 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6469 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6470 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6471 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6472 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6473 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6474 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6475 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6476 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6477 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6478 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6479 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6480 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6481 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6482 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6483 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6484 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6485 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6486 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6487 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6488 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6489 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6490 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6491 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6492 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6493 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6494 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6495 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6496 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6497 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6498 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6499 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6500 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6501 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6502 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6503 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6504 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6505 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6506 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6507 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6508 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6509 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6510 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6511 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6512 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6513 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6514 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6515 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6516 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6517 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6518 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6519 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6520 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6521 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6522 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6523 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6524 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6525 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6526 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6527 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6528 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6529 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6530 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6531 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6532 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6533 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6534 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6535 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6536 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6537 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6538 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6539 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6540 IREF ISBCS2 \$10007 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6541 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6542 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6543 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$6544 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$6545 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$6546 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$6547 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P PS=5.72U
+ PD=5.72U
M$6548 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6549 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P PS=3.62U
+ PD=2U
M$6550 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U
+ PD=3.62U
M$6551 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$6552 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6553 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6554 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6555 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6556 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6557 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6558 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6559 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6560 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6561 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6562 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6563 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6564 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6565 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6566 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6567 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6568 AVSS \$8587 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6569 \$7408 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6570 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6571 \$7673 \$8587 AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6572 AVSS \$8587 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6573 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6574 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6575 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6576 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6577 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6578 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6579 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6580 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6581 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6582 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6583 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6584 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6585 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6586 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6587 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6588 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6589 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6590 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6591 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6592 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6593 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6594 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6595 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6596 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6597 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6598 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6599 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6600 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6601 \$14873 \$9382 \$7673 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6602 \$7673 \$9382 \$14873 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6603 \$14873 \$9382 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6604 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6605 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6606 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6607 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6608 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6609 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6610 \$7408 \$9382 VOUT VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6611 VOUT \$9382 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6612 \$7408 \$9382 VOUT VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6613 \$14873 \$9382 \$7673 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6614 \$7673 \$9382 \$14873 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6615 \$14873 \$9382 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6616 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6617 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6618 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6619 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6620 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6621 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6622 VOUT \$9382 \$7408 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6623 \$7408 \$9382 VOUT VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6624 VOUT \$9382 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6625 \$14873 \$9382 \$7673 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6626 \$7673 \$9382 \$14873 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6627 \$14873 \$9382 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6628 \$7408 \$9382 VOUT VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6629 VOUT \$9382 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6630 \$7408 \$9382 VOUT VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6631 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6632 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6633 VOUT \$9382 \$7408 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6634 \$7408 \$9382 VOUT VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6635 VOUT \$9382 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6636 \$14873 \$9382 \$7673 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6637 \$7673 \$9382 \$14873 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6638 \$14873 \$9382 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6639 \$7408 \$9382 VOUT VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6640 VOUT \$9382 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6641 \$7408 \$9382 VOUT VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6642 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6643 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6644 \$14873 \$9382 \$7673 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6645 \$7673 \$9382 \$14873 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6646 \$14873 \$9382 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6647 VOUT \$9382 \$7408 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6648 \$7408 \$9382 VOUT VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6649 VOUT \$9382 \$7408 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6650 \$7673 \$9382 \$14873 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$6651 \$14873 \$9382 \$7673 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U
+ PD=2.8U
M$6652 \$7673 \$9382 \$14873 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$6653 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6654 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$6655 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6656 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6657 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6658 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6659 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6660 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6661 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$6662 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$6663 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6664 AVSS AVSS AVSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
C$6665 \$7674 \$7809 1.9208e-13 cap_mim_2f0_m4m5_noshield A=96.04P P=39.2U
C$6666 \$7675 \$7810 1.9208e-13 cap_mim_2f0_m4m5_noshield A=96.04P P=39.2U
C$6667 \$6456 \$6457 2e-11 cap_mim_2f0_m4m5_noshield A=10000P P=400U
C$6668 \$24406 \$24409 2e-11 cap_mim_2f0_m4m5_noshield A=10000P P=400U
.ENDS Filter_TOP
