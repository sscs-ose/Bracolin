* Extracted by KLayout with GF180MCU LVS runset on : 11/12/2023 13:14

.SUBCKT CM_n_net IN OUT8 OUT10 OUT12 OUT7 OUT9 OUT11 OUT2 OUT4 OUT6 OUT1 OUT3
+ OUT5 VSS
M$1 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$2 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$3 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$4 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$5 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$6 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$7 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$8 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$9 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$10 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$11 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$12 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$13 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$14 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$15 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$16 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$17 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$18 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$19 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$20 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$21 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$22 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$23 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$24 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$25 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$26 \$29 IN \$28 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$27 \$19 IN \$29 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$28 \$30 IN VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$29 \$31 IN \$30 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$30 \$32 IN \$19 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$31 \$33 IN \$32 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$32 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$33 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$34 \$35 IN \$34 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$35 \$20 IN \$35 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$36 \$36 IN VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$37 \$37 IN \$36 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$38 \$38 IN \$20 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$39 \$39 IN \$38 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$40 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$41 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$42 \$41 IN \$40 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$43 \$21 IN \$41 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$44 \$42 IN VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$45 \$43 IN \$42 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$46 \$44 IN \$21 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$47 \$45 IN \$44 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$48 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$49 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$50 \$64 IN \$28 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$51 \$65 IN \$64 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$52 \$67 IN \$66 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$53 \$31 IN \$67 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$54 \$69 IN \$68 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$55 \$33 IN \$69 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$56 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$57 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$58 \$70 IN \$34 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$59 \$71 IN \$70 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$60 \$73 IN \$72 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$61 \$37 IN \$73 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$62 \$75 IN \$74 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$63 \$39 IN \$75 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$64 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$65 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$66 \$76 IN \$40 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$67 \$77 IN \$76 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$68 \$79 IN \$78 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$69 \$43 IN \$79 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$70 \$81 IN \$80 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$71 \$45 IN \$81 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$72 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$73 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$74 \$110 IN \$109 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$75 \$65 IN \$110 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$76 \$111 IN \$66 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$77 \$100 IN \$111 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$78 \$112 IN \$68 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$79 \$113 IN \$112 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$80 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$81 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$82 \$115 IN \$114 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$83 \$71 IN \$115 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$84 \$116 IN \$72 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$85 \$101 IN \$116 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$86 \$117 IN \$74 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$87 \$118 IN \$117 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$88 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$89 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$90 \$120 IN \$119 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$91 \$77 IN \$120 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$92 \$121 IN \$78 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$93 \$102 IN \$121 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$94 \$122 IN \$80 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$95 \$123 IN \$122 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$96 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$97 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$98 \$151 IN \$109 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$99 \$152 IN \$151 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$100 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$101 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$102 \$154 IN \$153 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$103 \$113 IN \$154 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$104 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$105 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$106 \$155 IN \$114 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$107 \$156 IN \$155 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$108 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$109 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$110 \$158 IN \$157 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$111 \$118 IN \$158 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$112 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$113 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$114 \$159 IN \$119 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$115 \$160 IN \$159 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$116 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$117 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$118 \$162 IN \$161 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$119 \$123 IN \$162 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$120 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$121 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$122 \$191 IN OUT8 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$123 \$192 IN \$191 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$124 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$125 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$126 \$194 IN \$193 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$127 \$100 IN \$194 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$128 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$129 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$130 \$196 IN OUT10 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$131 \$197 IN \$196 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$132 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$133 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$134 \$199 IN \$198 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$135 \$101 IN \$199 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$136 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$137 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$138 \$201 IN OUT12 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$139 \$202 IN \$201 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$140 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$141 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$142 \$204 IN \$203 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$143 \$102 IN \$204 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$144 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$145 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$146 \$242 IN \$241 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$147 \$152 IN \$242 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$148 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$149 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$150 \$243 IN \$153 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$151 \$244 IN \$243 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$152 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$153 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$154 \$246 IN \$245 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$155 \$156 IN \$246 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$156 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$157 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$158 \$247 IN \$157 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$159 \$248 IN \$247 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$160 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$161 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$162 \$250 IN \$249 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$163 \$160 IN \$250 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$164 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$165 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$166 \$251 IN \$161 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$167 \$252 IN \$251 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$168 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$169 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$170 \$283 IN \$241 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$171 \$284 IN \$283 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$172 \$286 IN \$285 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$173 \$193 IN \$286 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$174 \$288 IN \$287 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$175 \$244 IN \$288 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$176 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$177 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$178 \$289 IN \$245 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$179 \$290 IN \$289 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$180 \$292 IN \$291 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$181 \$198 IN \$292 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$182 \$294 IN \$293 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$183 \$248 IN \$294 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$184 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$185 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$186 \$295 IN \$249 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$187 \$296 IN \$295 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$188 \$298 IN \$297 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$189 \$203 IN \$298 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$190 \$300 IN \$299 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$191 \$252 IN \$300 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$192 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$193 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$194 \$326 IN \$325 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$195 \$284 IN \$326 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$196 \$327 IN \$285 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$197 \$328 IN \$327 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$198 \$329 IN \$287 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$199 \$330 IN \$329 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$200 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$201 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$202 \$332 IN \$331 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$203 \$290 IN \$332 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$204 \$333 IN \$291 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$205 \$334 IN \$333 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$206 \$335 IN \$293 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$207 \$336 IN \$335 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$208 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$209 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$210 \$338 IN \$337 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$211 \$296 IN \$338 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$212 \$339 IN \$297 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$213 \$340 IN \$339 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$214 \$341 IN \$299 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$215 \$342 IN \$341 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$216 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$217 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$218 \$367 IN \$325 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$219 OUT7 IN \$367 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$220 \$369 IN \$192 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$221 \$328 IN \$369 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$222 \$370 IN VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$223 \$330 IN \$370 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$224 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$225 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$226 \$371 IN \$331 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$227 OUT9 IN \$371 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$228 \$373 IN \$197 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$229 \$334 IN \$373 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$230 \$374 IN VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$231 \$336 IN \$374 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$232 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$233 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$234 \$375 IN \$337 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$235 OUT11 IN \$375 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$236 \$377 IN \$202 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$237 \$340 IN \$377 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$238 \$378 IN VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$239 \$342 IN \$378 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$240 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$241 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$242 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$243 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$244 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$245 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$246 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$247 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$248 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$249 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$250 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$251 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$252 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$253 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$254 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$255 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$256 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$257 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$258 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$259 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$260 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$261 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$262 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$263 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$264 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$265 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$266 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$267 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$268 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$269 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$270 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$271 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$272 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$273 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$274 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$275 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$276 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$277 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$278 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$279 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$280 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$281 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$282 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$283 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$284 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$285 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$286 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$287 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$288 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$289 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$290 \$442 IN \$441 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$291 \$435 IN \$442 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$292 \$443 IN VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$293 \$444 IN \$443 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$294 \$445 IN \$435 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$295 \$446 IN \$445 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$296 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$297 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$298 \$448 IN \$447 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$299 \$436 IN \$448 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$300 \$449 IN VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$301 \$450 IN \$449 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$302 \$451 IN \$436 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$303 \$452 IN \$451 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$304 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$305 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$306 \$454 IN \$453 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$307 \$437 IN \$454 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$308 \$455 IN VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$309 \$456 IN \$455 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$310 \$457 IN \$437 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$311 \$458 IN \$457 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$312 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$313 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$314 \$480 IN \$441 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$315 \$481 IN \$480 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$316 \$483 IN \$482 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$317 \$444 IN \$483 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$318 \$485 IN \$484 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$319 \$446 IN \$485 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$320 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$321 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$322 \$486 IN \$447 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$323 \$487 IN \$486 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$324 \$489 IN \$488 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$325 \$450 IN \$489 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$326 \$491 IN \$490 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$327 \$452 IN \$491 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$328 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$329 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$330 \$492 IN \$453 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$331 \$493 IN \$492 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$332 \$495 IN \$494 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$333 \$456 IN \$495 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$334 \$497 IN \$496 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$335 \$458 IN \$497 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$336 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$337 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$338 \$526 IN \$525 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$339 \$481 IN \$526 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$340 \$527 IN \$482 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$341 \$516 IN \$527 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$342 \$528 IN \$484 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$343 \$529 IN \$528 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$344 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$345 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$346 \$531 IN \$530 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$347 \$487 IN \$531 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$348 \$532 IN \$488 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$349 \$517 IN \$532 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$350 \$533 IN \$490 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$351 \$534 IN \$533 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$352 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$353 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$354 \$536 IN \$535 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$355 \$493 IN \$536 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$356 \$537 IN \$494 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$357 \$518 IN \$537 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$358 \$538 IN \$496 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$359 \$539 IN \$538 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$360 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$361 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$362 \$567 IN \$525 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$363 \$568 IN \$567 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$364 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$365 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$366 \$570 IN \$569 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$367 \$529 IN \$570 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$368 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$369 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$370 \$571 IN \$530 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$371 \$572 IN \$571 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$372 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$373 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$374 \$574 IN \$573 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$375 \$534 IN \$574 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$376 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$377 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$378 \$575 IN \$535 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$379 \$576 IN \$575 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$380 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$381 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$382 \$578 IN \$577 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$383 \$539 IN \$578 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$384 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$385 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$386 \$607 IN OUT2 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$387 \$608 IN \$607 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$388 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$389 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$390 \$610 IN \$609 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$391 \$516 IN \$610 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$392 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$393 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$394 \$612 IN OUT4 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$395 \$613 IN \$612 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$396 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$397 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$398 \$615 IN \$614 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$399 \$517 IN \$615 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$400 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$401 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$402 \$617 IN OUT6 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$403 \$618 IN \$617 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$404 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$405 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$406 \$620 IN \$619 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$407 \$518 IN \$620 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$408 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$409 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$410 \$658 IN \$657 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$411 \$568 IN \$658 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$412 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$413 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$414 \$659 IN \$569 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$415 \$660 IN \$659 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$416 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$417 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$418 \$662 IN \$661 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$419 \$572 IN \$662 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$420 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$421 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$422 \$663 IN \$573 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$423 \$664 IN \$663 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$424 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$425 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$426 \$666 IN \$665 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$427 \$576 IN \$666 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$428 VSS IN IN VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$429 IN IN VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$430 \$667 IN \$577 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$431 \$668 IN \$667 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$432 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$433 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$434 \$699 IN \$657 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$435 \$700 IN \$699 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$436 \$702 IN \$701 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$437 \$609 IN \$702 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$438 \$704 IN \$703 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$439 \$660 IN \$704 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$440 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$441 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$442 \$705 IN \$661 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$443 \$706 IN \$705 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$444 \$708 IN \$707 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$445 \$614 IN \$708 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$446 \$710 IN \$709 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$447 \$664 IN \$710 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$448 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$449 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$450 \$711 IN \$665 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$451 \$712 IN \$711 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$452 \$714 IN \$713 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$453 \$619 IN \$714 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$454 \$716 IN \$715 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$455 \$668 IN \$716 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$456 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$457 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$458 \$742 IN \$741 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$459 \$700 IN \$742 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$460 \$743 IN \$701 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$461 \$744 IN \$743 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$462 \$745 IN \$703 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$463 \$746 IN \$745 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$464 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$465 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$466 \$748 IN \$747 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$467 \$706 IN \$748 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$468 \$749 IN \$707 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$469 \$750 IN \$749 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$470 \$751 IN \$709 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$471 \$752 IN \$751 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$472 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$473 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$474 \$754 IN \$753 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$475 \$712 IN \$754 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$476 \$755 IN \$713 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$477 \$756 IN \$755 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$478 \$757 IN \$715 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$479 \$758 IN \$757 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$480 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$481 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$482 \$783 IN \$741 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$483 OUT1 IN \$783 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$484 \$785 IN \$608 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$485 \$744 IN \$785 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$486 \$786 IN VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$487 \$746 IN \$786 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$488 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$489 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$490 \$787 IN \$747 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$491 OUT3 IN \$787 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$492 \$789 IN \$613 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$493 \$750 IN \$789 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$494 \$790 IN VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$495 \$752 IN \$790 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$496 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$497 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$498 \$791 IN \$753 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$499 OUT5 IN \$791 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$500 \$793 IN \$618 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$501 \$756 IN \$793 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$502 \$794 IN VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$503 \$758 IN \$794 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$504 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$505 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$506 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$507 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$508 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$509 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$510 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$511 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$512 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$513 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$514 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$515 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$516 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$517 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$518 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$519 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$520 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$521 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$522 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$523 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$524 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$525 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$526 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$527 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$528 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
.ENDS CM_n_net
