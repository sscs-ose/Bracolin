** sch_path: /home/gf180/Documents/gf180/gf180_work/PICO_contest/SAR_logic/xschem/D_reset_FF.sch
.subckt D_reset_FF VDDD VSSD Q nQ CLK D Reset Set
*.PININFO VDDD:B VSSD:B Q:B nQ:B CLK:I D:I Reset:I Set:I
x11 VDDD CLK nCLK VSSD inv_1x
x1 CLK_buf VDDD D net1 VSSD nCLK t_gate
x2 VDDD Set net2 net1 VSSD nor_2_1x
x4 nCLK VDDD net2 net4 VSSD CLK_buf t_gate
x6 VDDD Reset Q net4 VSSD nor_2_1x
x3 nCLK VDDD net3 net1 VSSD CLK_buf t_gate
x5 VDDD net2 net3 Reset VSSD nor_2_1x
x7 CLK_buf VDDD net5 net4 VSSD nCLK t_gate
x8 VDDD Q net5 Set VSSD nor_2_1x
x9 VDDD Q nQ VSSD inv_1x
x10 VDDD nCLK CLK_buf VSSD inv_1x
.ends

* expanding   symbol:  PICO_contest/SAR_logic/xschem/inv_1x.sym # of pins=4
** sym_path: /home/gf180/Documents/gf180/gf180_work/PICO_contest/SAR_logic/xschem/inv_1x.sym
** sch_path: /home/gf180/Documents/gf180/gf180_work/PICO_contest/SAR_logic/xschem/inv_1x.sch
.subckt inv_1x VDDD IN OUT VSSD
*.PININFO IN:I VDDD:B VSSD:B OUT:B
M1 OUT IN VDDD VDDD pfet_03v3 L=0.28u W=3.9u nf=1 m=1
M2 OUT IN VSSD VSSD nfet_03v3 L=0.28u W=1.56u nf=1 m=1
.ends


* expanding   symbol:  PICO_contest/SAR_logic/xschem/t_gate.sym # of pins=6
** sym_path: /home/gf180/Documents/gf180/gf180_work/PICO_contest/SAR_logic/xschem/t_gate.sym
** sch_path: /home/gf180/Documents/gf180/gf180_work/PICO_contest/SAR_logic/xschem/t_gate.sch
.subckt t_gate p_CLK VDDD IN OUT VSSD n_CLK
*.PININFO IN:B VDDD:B VSSD:B OUT:B n_CLK:I p_CLK:I
M1 IN n_CLK OUT VSSD nfet_03v3 L=0.28u W=1.56u nf=1 m=1
M2 IN p_CLK OUT VDDD pfet_03v3 L=0.28u W=3.9u nf=1 m=1
.ends


* expanding   symbol:  PICO_contest/SAR_logic/xschem/nor_2_1x.sym # of pins=5
** sym_path: /home/gf180/Documents/gf180/gf180_work/PICO_contest/SAR_logic/xschem/nor_2_1x.sym
** sch_path: /home/gf180/Documents/gf180/gf180_work/PICO_contest/SAR_logic/xschem/nor_2_1x.sch
.subckt nor_2_1x VDDD A OUT B VSSD
*.PININFO A:I B:I VDDD:B VSSD:B OUT:B
M1 OUT B VSSD VSSD nfet_03v3 L=0.28u W=1.56u nf=1 m=1
M2 OUT A VSSD VSSD nfet_03v3 L=0.28u W=1.56u nf=1 m=1
M3 OUT B net1 VDDD pfet_03v3 L=0.28u W=3.9u nf=1 m=1
M4 net1 A VDDD VDDD pfet_03v3 L=0.28u W=3.9u nf=1 m=1
.ends

.end
